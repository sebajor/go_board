// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jul 25 2020 17:39:27

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    o_Segment2_A,
    o_Segment1_E,
    o_UART_TX,
    o_Segment2_D,
    o_Segment1_F,
    o_Segment1_B,
    i_Clk,
    o_Segment2_G,
    o_Segment2_C,
    o_Segment1_G,
    o_Segment1_C,
    i_UART_RX,
    i_Switch_1,
    o_Segment2_F,
    o_Segment2_B,
    o_Segment1_D,
    o_LED_1,
    o_Segment2_E,
    o_Segment1_A);

    output o_Segment2_A;
    output o_Segment1_E;
    output o_UART_TX;
    output o_Segment2_D;
    output o_Segment1_F;
    output o_Segment1_B;
    input i_Clk;
    output o_Segment2_G;
    output o_Segment2_C;
    output o_Segment1_G;
    output o_Segment1_C;
    input i_UART_RX;
    input i_Switch_1;
    output o_Segment2_F;
    output o_Segment2_B;
    output o_Segment1_D;
    output o_LED_1;
    output o_Segment2_E;
    output o_Segment1_A;

    wire N__4755;
    wire N__4754;
    wire N__4753;
    wire N__4744;
    wire N__4743;
    wire N__4742;
    wire N__4735;
    wire N__4734;
    wire N__4733;
    wire N__4726;
    wire N__4725;
    wire N__4724;
    wire N__4717;
    wire N__4716;
    wire N__4715;
    wire N__4708;
    wire N__4707;
    wire N__4706;
    wire N__4699;
    wire N__4698;
    wire N__4697;
    wire N__4690;
    wire N__4689;
    wire N__4688;
    wire N__4681;
    wire N__4680;
    wire N__4679;
    wire N__4672;
    wire N__4671;
    wire N__4670;
    wire N__4663;
    wire N__4662;
    wire N__4661;
    wire N__4654;
    wire N__4653;
    wire N__4652;
    wire N__4645;
    wire N__4644;
    wire N__4643;
    wire N__4636;
    wire N__4635;
    wire N__4634;
    wire N__4627;
    wire N__4626;
    wire N__4625;
    wire N__4618;
    wire N__4617;
    wire N__4616;
    wire N__4609;
    wire N__4608;
    wire N__4607;
    wire N__4600;
    wire N__4599;
    wire N__4598;
    wire N__4591;
    wire N__4590;
    wire N__4589;
    wire N__4572;
    wire N__4571;
    wire N__4568;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4539;
    wire N__4536;
    wire N__4535;
    wire N__4532;
    wire N__4531;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4500;
    wire N__4497;
    wire N__4496;
    wire N__4495;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4464;
    wire N__4463;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4440;
    wire N__4437;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4406;
    wire N__4405;
    wire N__4402;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4380;
    wire N__4379;
    wire N__4378;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4366;
    wire N__4359;
    wire N__4358;
    wire N__4357;
    wire N__4356;
    wire N__4355;
    wire N__4354;
    wire N__4353;
    wire N__4352;
    wire N__4347;
    wire N__4346;
    wire N__4343;
    wire N__4338;
    wire N__4335;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4314;
    wire N__4305;
    wire N__4296;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4269;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4257;
    wire N__4256;
    wire N__4255;
    wire N__4254;
    wire N__4253;
    wire N__4252;
    wire N__4251;
    wire N__4250;
    wire N__4249;
    wire N__4248;
    wire N__4247;
    wire N__4246;
    wire N__4245;
    wire N__4244;
    wire N__4243;
    wire N__4242;
    wire N__4241;
    wire N__4240;
    wire N__4239;
    wire N__4238;
    wire N__4237;
    wire N__4236;
    wire N__4235;
    wire N__4234;
    wire N__4233;
    wire N__4232;
    wire N__4231;
    wire N__4230;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4154;
    wire N__4153;
    wire N__4152;
    wire N__4149;
    wire N__4142;
    wire N__4141;
    wire N__4140;
    wire N__4139;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4123;
    wire N__4116;
    wire N__4115;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4104;
    wire N__4103;
    wire N__4094;
    wire N__4093;
    wire N__4092;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4078;
    wire N__4071;
    wire N__4070;
    wire N__4069;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4055;
    wire N__4052;
    wire N__4045;
    wire N__4044;
    wire N__4043;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4024;
    wire N__4017;
    wire N__4014;
    wire N__4013;
    wire N__4012;
    wire N__4011;
    wire N__4008;
    wire N__4001;
    wire N__4000;
    wire N__3999;
    wire N__3998;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3982;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3948;
    wire N__3947;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3930;
    wire N__3929;
    wire N__3928;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3906;
    wire N__3903;
    wire N__3902;
    wire N__3901;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3879;
    wire N__3876;
    wire N__3875;
    wire N__3872;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3855;
    wire N__3852;
    wire N__3851;
    wire N__3850;
    wire N__3849;
    wire N__3846;
    wire N__3841;
    wire N__3838;
    wire N__3831;
    wire N__3828;
    wire N__3827;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3797;
    wire N__3796;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3784;
    wire N__3777;
    wire N__3774;
    wire N__3773;
    wire N__3772;
    wire N__3769;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3747;
    wire N__3744;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3659;
    wire N__3656;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3621;
    wire N__3618;
    wire N__3617;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3578;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3564;
    wire N__3561;
    wire N__3560;
    wire N__3559;
    wire N__3558;
    wire N__3555;
    wire N__3548;
    wire N__3543;
    wire N__3540;
    wire N__3539;
    wire N__3538;
    wire N__3537;
    wire N__3528;
    wire N__3527;
    wire N__3526;
    wire N__3525;
    wire N__3522;
    wire N__3521;
    wire N__3520;
    wire N__3513;
    wire N__3510;
    wire N__3507;
    wire N__3504;
    wire N__3503;
    wire N__3500;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3488;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3471;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3452;
    wire N__3447;
    wire N__3446;
    wire N__3445;
    wire N__3442;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3426;
    wire N__3425;
    wire N__3422;
    wire N__3421;
    wire N__3420;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3412;
    wire N__3411;
    wire N__3410;
    wire N__3409;
    wire N__3408;
    wire N__3401;
    wire N__3396;
    wire N__3385;
    wire N__3378;
    wire N__3375;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3363;
    wire N__3362;
    wire N__3361;
    wire N__3360;
    wire N__3359;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3338;
    wire N__3327;
    wire N__3326;
    wire N__3325;
    wire N__3324;
    wire N__3323;
    wire N__3322;
    wire N__3321;
    wire N__3318;
    wire N__3311;
    wire N__3304;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3245;
    wire N__3244;
    wire N__3243;
    wire N__3240;
    wire N__3233;
    wire N__3232;
    wire N__3231;
    wire N__3230;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3201;
    wire N__3198;
    wire N__3197;
    wire N__3196;
    wire N__3195;
    wire N__3192;
    wire N__3185;
    wire N__3184;
    wire N__3183;
    wire N__3182;
    wire N__3181;
    wire N__3178;
    wire N__3175;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3153;
    wire N__3152;
    wire N__3151;
    wire N__3148;
    wire N__3147;
    wire N__3146;
    wire N__3143;
    wire N__3142;
    wire N__3141;
    wire N__3138;
    wire N__3137;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3099;
    wire N__3098;
    wire N__3097;
    wire N__3096;
    wire N__3095;
    wire N__3094;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3077;
    wire N__3074;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3012;
    wire N__3009;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2945;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2904;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2894;
    wire N__2893;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2881;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2867;
    wire N__2864;
    wire N__2861;
    wire N__2856;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2835;
    wire N__2834;
    wire N__2829;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2817;
    wire N__2816;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2806;
    wire N__2805;
    wire N__2802;
    wire N__2797;
    wire N__2794;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2769;
    wire N__2766;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2754;
    wire N__2751;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2739;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2721;
    wire N__2720;
    wire N__2717;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2700;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2685;
    wire N__2684;
    wire N__2683;
    wire N__2680;
    wire N__2675;
    wire N__2670;
    wire N__2669;
    wire N__2668;
    wire N__2665;
    wire N__2660;
    wire N__2655;
    wire N__2652;
    wire N__2651;
    wire N__2650;
    wire N__2649;
    wire N__2646;
    wire N__2643;
    wire N__2638;
    wire N__2631;
    wire N__2628;
    wire N__2627;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2610;
    wire N__2607;
    wire N__2606;
    wire N__2605;
    wire N__2604;
    wire N__2603;
    wire N__2600;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2580;
    wire N__2577;
    wire N__2576;
    wire N__2575;
    wire N__2574;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2544;
    wire N__2541;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2529;
    wire N__2526;
    wire N__2525;
    wire N__2524;
    wire N__2523;
    wire N__2520;
    wire N__2517;
    wire N__2514;
    wire N__2511;
    wire N__2502;
    wire N__2501;
    wire N__2500;
    wire N__2499;
    wire N__2496;
    wire N__2493;
    wire N__2490;
    wire N__2487;
    wire N__2478;
    wire N__2475;
    wire N__2474;
    wire N__2469;
    wire N__2466;
    wire N__2465;
    wire N__2464;
    wire N__2463;
    wire N__2462;
    wire N__2461;
    wire N__2458;
    wire N__2455;
    wire N__2452;
    wire N__2445;
    wire N__2442;
    wire N__2433;
    wire N__2432;
    wire N__2431;
    wire N__2430;
    wire N__2429;
    wire N__2428;
    wire N__2425;
    wire N__2418;
    wire N__2415;
    wire N__2412;
    wire N__2403;
    wire N__2402;
    wire N__2397;
    wire N__2394;
    wire N__2393;
    wire N__2392;
    wire N__2391;
    wire N__2390;
    wire N__2389;
    wire N__2388;
    wire N__2383;
    wire N__2380;
    wire N__2379;
    wire N__2378;
    wire N__2375;
    wire N__2368;
    wire N__2363;
    wire N__2358;
    wire N__2349;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2337;
    wire N__2336;
    wire N__2335;
    wire N__2334;
    wire N__2331;
    wire N__2326;
    wire N__2323;
    wire N__2316;
    wire N__2315;
    wire N__2314;
    wire N__2313;
    wire N__2312;
    wire N__2309;
    wire N__2308;
    wire N__2305;
    wire N__2304;
    wire N__2303;
    wire N__2302;
    wire N__2299;
    wire N__2292;
    wire N__2287;
    wire N__2284;
    wire N__2281;
    wire N__2278;
    wire N__2277;
    wire N__2270;
    wire N__2267;
    wire N__2262;
    wire N__2259;
    wire N__2258;
    wire N__2251;
    wire N__2246;
    wire N__2241;
    wire N__2238;
    wire N__2235;
    wire N__2232;
    wire N__2229;
    wire N__2226;
    wire N__2223;
    wire N__2220;
    wire N__2219;
    wire N__2216;
    wire N__2213;
    wire N__2212;
    wire N__2207;
    wire N__2204;
    wire N__2199;
    wire N__2196;
    wire N__2193;
    wire N__2190;
    wire N__2187;
    wire N__2184;
    wire N__2181;
    wire N__2178;
    wire N__2175;
    wire N__2172;
    wire N__2169;
    wire N__2166;
    wire N__2163;
    wire N__2160;
    wire N__2157;
    wire N__2156;
    wire N__2153;
    wire N__2150;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2136;
    wire N__2133;
    wire N__2132;
    wire N__2129;
    wire N__2126;
    wire N__2121;
    wire N__2118;
    wire N__2115;
    wire N__2114;
    wire N__2113;
    wire N__2108;
    wire N__2105;
    wire N__2100;
    wire N__2097;
    wire N__2094;
    wire N__2093;
    wire N__2088;
    wire N__2085;
    wire N__2082;
    wire N__2079;
    wire N__2076;
    wire N__2073;
    wire N__2070;
    wire N__2067;
    wire N__2066;
    wire N__2065;
    wire N__2060;
    wire N__2057;
    wire N__2052;
    wire N__2051;
    wire N__2050;
    wire N__2049;
    wire N__2042;
    wire N__2039;
    wire N__2034;
    wire N__2031;
    wire N__2028;
    wire N__2025;
    wire N__2024;
    wire N__2019;
    wire N__2018;
    wire N__2015;
    wire N__2012;
    wire N__2007;
    wire N__2004;
    wire N__2003;
    wire N__1998;
    wire N__1995;
    wire N__1992;
    wire N__1991;
    wire N__1990;
    wire N__1987;
    wire N__1984;
    wire N__1983;
    wire N__1980;
    wire N__1977;
    wire N__1974;
    wire N__1971;
    wire N__1962;
    wire N__1959;
    wire N__1958;
    wire N__1957;
    wire N__1956;
    wire N__1951;
    wire N__1946;
    wire N__1941;
    wire N__1938;
    wire N__1937;
    wire N__1932;
    wire N__1929;
    wire N__1926;
    wire N__1923;
    wire N__1920;
    wire N__1917;
    wire N__1914;
    wire N__1911;
    wire N__1908;
    wire N__1905;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_10_0_;
    wire \uart_rx.un1_index_cry_0 ;
    wire \uart_rx.un1_index_cry_1 ;
    wire \uart_rx.un1_index_cry_2 ;
    wire \uart_rx.r_datace_0_2 ;
    wire \uart_rx.N_146_cascade_ ;
    wire \uart_rx.N_146 ;
    wire \uart_rx.state_srsts_i_a2_3_3_cascade_ ;
    wire \uart_rx.state_srsts_0_a2_2_4 ;
    wire \uart_rx.N_147_cascade_ ;
    wire \uart_rx.state_srsts_0_a2_1_4 ;
    wire \uart_rx.N_136_cascade_ ;
    wire \uart_rx.stateZ0Z_5 ;
    wire \uart_rx.state_srsts_0_a2_0_2_2_cascade_ ;
    wire \uart_rx.stateZ0Z_3 ;
    wire \uart_rx.N_136 ;
    wire \uart_rx.state_nss_0_i_1_0 ;
    wire \uart_rx.state_srsts_i_o2_1_1 ;
    wire \uart_rx.state_srsts_i_a2_1_0_1_cascade_ ;
    wire \uart_rx.state_srsts_0_a2_0_1_0_2 ;
    wire \uart_rx.N_130_cascade_ ;
    wire \uart_rx.N_109_0 ;
    wire \uart_rx.stateZ0Z_1 ;
    wire \uart_rx.state_srsts_0_a2_0_1_4 ;
    wire \uart_rx.state_srsts_0_a2_0_1_4_cascade_ ;
    wire \uart_rx.timer_RNIUELTZ0Z_0 ;
    wire r_disp2_i_1;
    wire r_disp2_i_0;
    wire r_disp2_i_6;
    wire r_disp2_i_5;
    wire r_disp1_i_1;
    wire \uart_rx.r_dataZ1Z_2 ;
    wire \uart_rx.r_dataZ1Z_0 ;
    wire r_disp1_i_6;
    wire \uart_rx.N_139 ;
    wire \uart_rx.indexZ0Z_3 ;
    wire \uart_rx.indexZ0Z_1 ;
    wire \uart_rx.r_datace_0_6 ;
    wire \uart_rx.indexZ0Z_2 ;
    wire \uart_rx.indexZ0Z_0 ;
    wire \uart_rx.r_datace_0_3 ;
    wire \uart_rx.N_122_i ;
    wire \uart_rx.N_147 ;
    wire \uart_rx.N_142 ;
    wire i_UART_RX_c;
    wire \uart_rx.r_datace_0_5 ;
    wire \uart_rx.state_isoZ0Z_0 ;
    wire \uart_rx.stateZ0Z_2 ;
    wire \uart_rx.N_123_i ;
    wire \uart_rx.timerZ0Z_0 ;
    wire bfn_2_12_0_;
    wire \uart_rx.timerZ0Z_1 ;
    wire \uart_rx.un1_timer_cry_0 ;
    wire \uart_rx.timerZ0Z_2 ;
    wire \uart_rx.un1_timer_cry_1 ;
    wire \uart_rx.timerZ0Z_3 ;
    wire \uart_rx.un1_timer_cry_2 ;
    wire \uart_rx.timerZ0Z_4 ;
    wire \uart_rx.un1_timer_cry_3 ;
    wire \uart_rx.timerZ0Z_5 ;
    wire \uart_rx.un1_timer_cry_4 ;
    wire \uart_rx.timerZ0Z_6 ;
    wire \uart_rx.un1_timer_cry_5 ;
    wire \uart_rx.timerZ0Z_7 ;
    wire \uart_rx.un1_timer_cry_6 ;
    wire \uart_rx.un1_timer_cry_7 ;
    wire bfn_2_13_0_;
    wire \uart_rx.timerZ0Z_8 ;
    wire \uart_rx.state_RNIQRIGZ0Z_2 ;
    wire \uart_rx.stateZ0Z_6 ;
    wire \uart_rx.stateZ0Z_0 ;
    wire \uart_rx.r_dataZ0Z_7 ;
    wire \uart_rx.r_dataZ0Z_6 ;
    wire \uart_rx.r_dataZ1Z_1 ;
    wire \uart_rx.r_dataZ0Z_3 ;
    wire \uart_rx.r_dataZ0Z_4 ;
    wire r_disp1_i_5;
    wire r_disp1_i_4;
    wire CONSTANT_ONE_NET;
    wire \uart_tx.r_dataZ0Z_8 ;
    wire \uart_tx.r_dataZ0Z_0 ;
    wire \uart_tx.r_dataZ0Z_5 ;
    wire \uart_tx.out_data_2_4_i_m2_ns_1_cascade_ ;
    wire \uart_tx.r_dataZ0Z_1 ;
    wire \uart_tx.r_dataZ0Z_4 ;
    wire r_uart_charZ0Z_0;
    wire r_uart_charZ0Z_1;
    wire r_uart_charZ0Z_4;
    wire r_uart_charZ0Z_5;
    wire valid_msg_0;
    wire r_disp1_i_0;
    wire r_disp1_i_3;
    wire uart_data_0;
    wire uart_data_2;
    wire uart_data_1;
    wire uart_data_3;
    wire r_disp1_i_2;
    wire \uart_tx.counter12_6_0_cascade_ ;
    wire \uart_tx.g0_rn_0 ;
    wire \uart_tx.g0_sn ;
    wire \uart_tx.next_state_1_0_m2_i_a2_1_3_0 ;
    wire \uart_tx.next_state_1_0_m2_i_0_0_cascade_ ;
    wire \uart_tx.g0_0_3 ;
    wire \uart_tx.counter12_7_3_cascade_ ;
    wire \uart_tx.counter12_7 ;
    wire \uart_tx.counter12_7_cascade_ ;
    wire valid_msg;
    wire o_LED_1_c;
    wire uart_rx_tvalidZ0;
    wire \uart_tx.stateZ0Z_0 ;
    wire \uart_tx.un1_index_ac0_1_0 ;
    wire \uart_tx.indexZ0Z_2 ;
    wire \uart_tx.indexZ0Z_0 ;
    wire \uart_tx.out_data_2_5_i_m2_ns_1_cascade_ ;
    wire \uart_tx.N_57 ;
    wire \uart_tx.indexZ0Z_1 ;
    wire \uart_tx.N_56_cascade_ ;
    wire \uart_tx.indexZ0Z_3 ;
    wire \uart_tx.N_55_cascade_ ;
    wire \uart_tx.out_data_3_iv_0_a2_1 ;
    wire o_UART_TX_c;
    wire r_uart_charZ0Z_2;
    wire \uart_tx.r_dataZ0Z_2 ;
    wire r_uart_charZ0Z_3;
    wire \uart_tx.r_dataZ0Z_3 ;
    wire r_uart_charZ0Z_6;
    wire \uart_tx.r_dataZ0Z_6 ;
    wire r_uart_charZ0Z_7;
    wire \uart_tx.r_dataZ0Z_7 ;
    wire \uart_tx.r_data_0_sqmuxa ;
    wire \uart_rx.r_dataZ0Z_5 ;
    wire \uart_rx.state_RNIIKQGZ0Z_6 ;
    wire r_disp2_i_2;
    wire r_disp2_i_3;
    wire uart_data_6;
    wire uart_data_5;
    wire uart_data_7;
    wire uart_data_4;
    wire r_disp2_i_4;
    wire \uart_tx.N_50 ;
    wire \uart_tx.counterZ0Z_0 ;
    wire bfn_6_9_0_;
    wire \uart_tx.counterZ0Z_1 ;
    wire \uart_tx.un1_counter_5_cry_0 ;
    wire \uart_tx.counterZ0Z_2 ;
    wire \uart_tx.un1_counter_5_cry_1 ;
    wire \uart_tx.counterZ0Z_3 ;
    wire \uart_tx.un1_counter_5_cry_2 ;
    wire \uart_tx.counterZ0Z_4 ;
    wire \uart_tx.un1_counter_5_cry_3 ;
    wire \uart_tx.counterZ0Z_5 ;
    wire \uart_tx.un1_counter_5_cry_4 ;
    wire \uart_tx.counterZ0Z_6 ;
    wire \uart_tx.un1_counter_5_cry_5 ;
    wire \uart_tx.counterZ0Z_7 ;
    wire \uart_tx.un1_counter_5_cry_6 ;
    wire \uart_tx.un1_counter_5_cry_7 ;
    wire \uart_tx.counterZ0Z_8 ;
    wire bfn_6_10_0_;
    wire \uart_tx.un1_counter_5_cry_8 ;
    wire \uart_tx.counterZ0Z_9 ;
    wire \uart_tx.state_RNICAH01Z0Z_0 ;
    wire \uart_tx.counter_RNI6M34Z0Z_1 ;
    wire \uart_tx.counter_RNI1V9O_0Z0Z_4 ;
    wire \uart_tx.counter12_6 ;
    wire \uart_tx.N_29 ;
    wire \uart_tx.stateZ0Z_1 ;
    wire \uart_tx.tready5 ;
    wire uart_tx_tready;
    wire i_Clk_c_g;
    wire _gnd_net_;

    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__4753),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__4755),
            .DIN(N__4754),
            .DOUT(N__4753),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__4755),
            .PADOUT(N__4754),
            .PADIN(N__4753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_F_obuf_iopad (
            .OE(N__4744),
            .DIN(N__4743),
            .DOUT(N__4742),
            .PACKAGEPIN(o_Segment2_F));
    defparam o_Segment2_F_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_F_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_F_obuf_preio (
            .PADOEN(N__4744),
            .PADOUT(N__4743),
            .PADIN(N__4742),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2169),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_1_obuf_iopad (
            .OE(N__4735),
            .DIN(N__4734),
            .DOUT(N__4733),
            .PACKAGEPIN(o_LED_1));
    defparam o_LED_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_1_obuf_preio (
            .PADOEN(N__4735),
            .PADOUT(N__4734),
            .PADIN(N__4733),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3471),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_B_obuf_iopad (
            .OE(N__4726),
            .DIN(N__4725),
            .DOUT(N__4724),
            .PACKAGEPIN(o_Segment2_B));
    defparam o_Segment2_B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_B_obuf_preio (
            .PADOEN(N__4726),
            .PADOUT(N__4725),
            .PADIN(N__4724),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2940),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_G_obuf_iopad (
            .OE(N__4717),
            .DIN(N__4716),
            .DOUT(N__4715),
            .PACKAGEPIN(o_Segment1_G));
    defparam o_Segment1_G_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_G_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_G_obuf_preio (
            .PADOEN(N__4717),
            .PADOUT(N__4716),
            .PADIN(N__4715),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_C_obuf_iopad (
            .OE(N__4708),
            .DIN(N__4707),
            .DOUT(N__4706),
            .PACKAGEPIN(o_Segment1_C));
    defparam o_Segment1_C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_C_obuf_preio (
            .PADOEN(N__4708),
            .PADOUT(N__4707),
            .PADIN(N__4706),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3975),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_1_ibuf_iopad (
            .OE(N__4699),
            .DIN(N__4698),
            .DOUT(N__4697),
            .PACKAGEPIN(i_Switch_1));
    defparam i_Switch_1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_1_ibuf_preio (
            .PADOEN(N__4699),
            .PADOUT(N__4698),
            .PADIN(N__4697),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(o_LED_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_B_obuf_iopad (
            .OE(N__4690),
            .DIN(N__4689),
            .DOUT(N__4688),
            .PACKAGEPIN(o_Segment1_B));
    defparam o_Segment1_B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_B_obuf_preio (
            .PADOEN(N__4690),
            .PADOUT(N__4689),
            .PADIN(N__4688),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2175),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_D_obuf_iopad (
            .OE(N__4681),
            .DIN(N__4680),
            .DOUT(N__4679),
            .PACKAGEPIN(o_Segment1_D));
    defparam o_Segment1_D_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_D_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_D_obuf_preio (
            .PADOEN(N__4681),
            .PADOUT(N__4680),
            .PADIN(N__4679),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4167),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_F_obuf_iopad (
            .OE(N__4672),
            .DIN(N__4671),
            .DOUT(N__4670),
            .PACKAGEPIN(o_Segment1_F));
    defparam o_Segment1_F_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_F_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_F_obuf_preio (
            .PADOEN(N__4672),
            .PADOUT(N__4671),
            .PADIN(N__4670),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2193),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_E_obuf_iopad (
            .OE(N__4663),
            .DIN(N__4662),
            .DOUT(N__4661),
            .PACKAGEPIN(o_Segment1_E));
    defparam o_Segment1_E_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_E_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_E_obuf_preio (
            .PADOEN(N__4663),
            .PADOUT(N__4662),
            .PADIN(N__4661),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3594),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_A_obuf_iopad (
            .OE(N__4654),
            .DIN(N__4653),
            .DOUT(N__4652),
            .PACKAGEPIN(o_Segment2_A));
    defparam o_Segment2_A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_A_obuf_preio (
            .PADOEN(N__4654),
            .PADOUT(N__4653),
            .PADIN(N__4652),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2121),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_G_obuf_iopad (
            .OE(N__4645),
            .DIN(N__4644),
            .DOUT(N__4643),
            .PACKAGEPIN(o_Segment2_G));
    defparam o_Segment2_G_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_G_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_G_obuf_preio (
            .PADOEN(N__4645),
            .PADOUT(N__4644),
            .PADIN(N__4643),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3267),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_D_obuf_iopad (
            .OE(N__4636),
            .DIN(N__4635),
            .DOUT(N__4634),
            .PACKAGEPIN(o_Segment2_D));
    defparam o_Segment2_D_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_D_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_D_obuf_preio (
            .PADOEN(N__4636),
            .PADOUT(N__4635),
            .PADIN(N__4634),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_UART_TX_obuf_iopad (
            .OE(N__4627),
            .DIN(N__4626),
            .DOUT(N__4625),
            .PACKAGEPIN(o_UART_TX));
    defparam o_UART_TX_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_UART_TX_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_UART_TX_obuf_preio (
            .PADOEN(N__4627),
            .PADOUT(N__4626),
            .PADIN(N__4625),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3732),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_E_obuf_iopad (
            .OE(N__4618),
            .DIN(N__4617),
            .DOUT(N__4616),
            .PACKAGEPIN(o_Segment2_E));
    defparam o_Segment2_E_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_E_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_E_obuf_preio (
            .PADOEN(N__4618),
            .PADOUT(N__4617),
            .PADIN(N__4616),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3036),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_C_obuf_iopad (
            .OE(N__4609),
            .DIN(N__4608),
            .DOUT(N__4607),
            .PACKAGEPIN(o_Segment2_C));
    defparam o_Segment2_C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_C_obuf_preio (
            .PADOEN(N__4609),
            .PADOUT(N__4608),
            .PADIN(N__4607),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2934),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_UART_RX_ibuf_iopad (
            .OE(N__4600),
            .DIN(N__4599),
            .DOUT(N__4598),
            .PACKAGEPIN(i_UART_RX));
    defparam i_UART_RX_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_UART_RX_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_UART_RX_ibuf_preio (
            .PADOEN(N__4600),
            .PADOUT(N__4599),
            .PADIN(N__4598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_UART_RX_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_A_obuf_iopad (
            .OE(N__4591),
            .DIN(N__4590),
            .DOUT(N__4589),
            .PACKAGEPIN(o_Segment1_A));
    defparam o_Segment1_A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_A_obuf_preio (
            .PADOEN(N__4591),
            .PADOUT(N__4590),
            .PADIN(N__4589),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2181),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1053 (
            .O(N__4572),
            .I(N__4568));
    CascadeMux I__1052 (
            .O(N__4571),
            .I(N__4564));
    LocalMux I__1051 (
            .O(N__4568),
            .I(N__4561));
    InMux I__1050 (
            .O(N__4567),
            .I(N__4557));
    InMux I__1049 (
            .O(N__4564),
            .I(N__4554));
    Span4Mux_h I__1048 (
            .O(N__4561),
            .I(N__4551));
    InMux I__1047 (
            .O(N__4560),
            .I(N__4548));
    LocalMux I__1046 (
            .O(N__4557),
            .I(\uart_tx.counterZ0Z_6 ));
    LocalMux I__1045 (
            .O(N__4554),
            .I(\uart_tx.counterZ0Z_6 ));
    Odrv4 I__1044 (
            .O(N__4551),
            .I(\uart_tx.counterZ0Z_6 ));
    LocalMux I__1043 (
            .O(N__4548),
            .I(\uart_tx.counterZ0Z_6 ));
    InMux I__1042 (
            .O(N__4539),
            .I(\uart_tx.un1_counter_5_cry_5 ));
    CascadeMux I__1041 (
            .O(N__4536),
            .I(N__4532));
    CascadeMux I__1040 (
            .O(N__4535),
            .I(N__4527));
    InMux I__1039 (
            .O(N__4532),
            .I(N__4524));
    CascadeMux I__1038 (
            .O(N__4531),
            .I(N__4521));
    InMux I__1037 (
            .O(N__4530),
            .I(N__4518));
    InMux I__1036 (
            .O(N__4527),
            .I(N__4515));
    LocalMux I__1035 (
            .O(N__4524),
            .I(N__4512));
    InMux I__1034 (
            .O(N__4521),
            .I(N__4509));
    LocalMux I__1033 (
            .O(N__4518),
            .I(\uart_tx.counterZ0Z_7 ));
    LocalMux I__1032 (
            .O(N__4515),
            .I(\uart_tx.counterZ0Z_7 ));
    Odrv4 I__1031 (
            .O(N__4512),
            .I(\uart_tx.counterZ0Z_7 ));
    LocalMux I__1030 (
            .O(N__4509),
            .I(\uart_tx.counterZ0Z_7 ));
    InMux I__1029 (
            .O(N__4500),
            .I(\uart_tx.un1_counter_5_cry_6 ));
    InMux I__1028 (
            .O(N__4497),
            .I(N__4491));
    InMux I__1027 (
            .O(N__4496),
            .I(N__4488));
    InMux I__1026 (
            .O(N__4495),
            .I(N__4485));
    InMux I__1025 (
            .O(N__4494),
            .I(N__4482));
    LocalMux I__1024 (
            .O(N__4491),
            .I(\uart_tx.counterZ0Z_8 ));
    LocalMux I__1023 (
            .O(N__4488),
            .I(\uart_tx.counterZ0Z_8 ));
    LocalMux I__1022 (
            .O(N__4485),
            .I(\uart_tx.counterZ0Z_8 ));
    LocalMux I__1021 (
            .O(N__4482),
            .I(\uart_tx.counterZ0Z_8 ));
    InMux I__1020 (
            .O(N__4473),
            .I(bfn_6_10_0_));
    InMux I__1019 (
            .O(N__4470),
            .I(\uart_tx.un1_counter_5_cry_8 ));
    CascadeMux I__1018 (
            .O(N__4467),
            .I(N__4464));
    InMux I__1017 (
            .O(N__4464),
            .I(N__4459));
    CascadeMux I__1016 (
            .O(N__4463),
            .I(N__4456));
    InMux I__1015 (
            .O(N__4462),
            .I(N__4453));
    LocalMux I__1014 (
            .O(N__4459),
            .I(N__4450));
    InMux I__1013 (
            .O(N__4456),
            .I(N__4447));
    LocalMux I__1012 (
            .O(N__4453),
            .I(\uart_tx.counterZ0Z_9 ));
    Odrv4 I__1011 (
            .O(N__4450),
            .I(\uart_tx.counterZ0Z_9 ));
    LocalMux I__1010 (
            .O(N__4447),
            .I(\uart_tx.counterZ0Z_9 ));
    SRMux I__1009 (
            .O(N__4440),
            .I(N__4437));
    LocalMux I__1008 (
            .O(N__4437),
            .I(N__4433));
    SRMux I__1007 (
            .O(N__4436),
            .I(N__4430));
    Span4Mux_v I__1006 (
            .O(N__4433),
            .I(N__4425));
    LocalMux I__1005 (
            .O(N__4430),
            .I(N__4425));
    Odrv4 I__1004 (
            .O(N__4425),
            .I(\uart_tx.state_RNICAH01Z0Z_0 ));
    InMux I__1003 (
            .O(N__4422),
            .I(N__4419));
    LocalMux I__1002 (
            .O(N__4419),
            .I(\uart_tx.counter_RNI6M34Z0Z_1 ));
    CascadeMux I__1001 (
            .O(N__4416),
            .I(N__4413));
    InMux I__1000 (
            .O(N__4413),
            .I(N__4410));
    LocalMux I__999 (
            .O(N__4410),
            .I(\uart_tx.counter_RNI1V9O_0Z0Z_4 ));
    InMux I__998 (
            .O(N__4407),
            .I(N__4402));
    InMux I__997 (
            .O(N__4406),
            .I(N__4398));
    InMux I__996 (
            .O(N__4405),
            .I(N__4395));
    LocalMux I__995 (
            .O(N__4402),
            .I(N__4392));
    InMux I__994 (
            .O(N__4401),
            .I(N__4389));
    LocalMux I__993 (
            .O(N__4398),
            .I(\uart_tx.counter12_6 ));
    LocalMux I__992 (
            .O(N__4395),
            .I(\uart_tx.counter12_6 ));
    Odrv4 I__991 (
            .O(N__4392),
            .I(\uart_tx.counter12_6 ));
    LocalMux I__990 (
            .O(N__4389),
            .I(\uart_tx.counter12_6 ));
    InMux I__989 (
            .O(N__4380),
            .I(N__4374));
    InMux I__988 (
            .O(N__4379),
            .I(N__4371));
    InMux I__987 (
            .O(N__4378),
            .I(N__4366));
    InMux I__986 (
            .O(N__4377),
            .I(N__4366));
    LocalMux I__985 (
            .O(N__4374),
            .I(\uart_tx.N_29 ));
    LocalMux I__984 (
            .O(N__4371),
            .I(\uart_tx.N_29 ));
    LocalMux I__983 (
            .O(N__4366),
            .I(\uart_tx.N_29 ));
    InMux I__982 (
            .O(N__4359),
            .I(N__4347));
    InMux I__981 (
            .O(N__4358),
            .I(N__4347));
    InMux I__980 (
            .O(N__4357),
            .I(N__4343));
    InMux I__979 (
            .O(N__4356),
            .I(N__4338));
    InMux I__978 (
            .O(N__4355),
            .I(N__4338));
    InMux I__977 (
            .O(N__4354),
            .I(N__4335));
    CascadeMux I__976 (
            .O(N__4353),
            .I(N__4331));
    CascadeMux I__975 (
            .O(N__4352),
            .I(N__4328));
    LocalMux I__974 (
            .O(N__4347),
            .I(N__4324));
    InMux I__973 (
            .O(N__4346),
            .I(N__4321));
    LocalMux I__972 (
            .O(N__4343),
            .I(N__4314));
    LocalMux I__971 (
            .O(N__4338),
            .I(N__4314));
    LocalMux I__970 (
            .O(N__4335),
            .I(N__4314));
    InMux I__969 (
            .O(N__4334),
            .I(N__4305));
    InMux I__968 (
            .O(N__4331),
            .I(N__4305));
    InMux I__967 (
            .O(N__4328),
            .I(N__4305));
    InMux I__966 (
            .O(N__4327),
            .I(N__4305));
    Odrv4 I__965 (
            .O(N__4324),
            .I(\uart_tx.stateZ0Z_1 ));
    LocalMux I__964 (
            .O(N__4321),
            .I(\uart_tx.stateZ0Z_1 ));
    Odrv4 I__963 (
            .O(N__4314),
            .I(\uart_tx.stateZ0Z_1 ));
    LocalMux I__962 (
            .O(N__4305),
            .I(\uart_tx.stateZ0Z_1 ));
    SRMux I__961 (
            .O(N__4296),
            .I(N__4292));
    SRMux I__960 (
            .O(N__4295),
            .I(N__4289));
    LocalMux I__959 (
            .O(N__4292),
            .I(N__4286));
    LocalMux I__958 (
            .O(N__4289),
            .I(N__4282));
    Span4Mux_h I__957 (
            .O(N__4286),
            .I(N__4279));
    InMux I__956 (
            .O(N__4285),
            .I(N__4276));
    Odrv4 I__955 (
            .O(N__4282),
            .I(\uart_tx.tready5 ));
    Odrv4 I__954 (
            .O(N__4279),
            .I(\uart_tx.tready5 ));
    LocalMux I__953 (
            .O(N__4276),
            .I(\uart_tx.tready5 ));
    InMux I__952 (
            .O(N__4269),
            .I(N__4265));
    InMux I__951 (
            .O(N__4268),
            .I(N__4262));
    LocalMux I__950 (
            .O(N__4265),
            .I(uart_tx_tready));
    LocalMux I__949 (
            .O(N__4262),
            .I(uart_tx_tready));
    ClkMux I__948 (
            .O(N__4257),
            .I(N__4173));
    ClkMux I__947 (
            .O(N__4256),
            .I(N__4173));
    ClkMux I__946 (
            .O(N__4255),
            .I(N__4173));
    ClkMux I__945 (
            .O(N__4254),
            .I(N__4173));
    ClkMux I__944 (
            .O(N__4253),
            .I(N__4173));
    ClkMux I__943 (
            .O(N__4252),
            .I(N__4173));
    ClkMux I__942 (
            .O(N__4251),
            .I(N__4173));
    ClkMux I__941 (
            .O(N__4250),
            .I(N__4173));
    ClkMux I__940 (
            .O(N__4249),
            .I(N__4173));
    ClkMux I__939 (
            .O(N__4248),
            .I(N__4173));
    ClkMux I__938 (
            .O(N__4247),
            .I(N__4173));
    ClkMux I__937 (
            .O(N__4246),
            .I(N__4173));
    ClkMux I__936 (
            .O(N__4245),
            .I(N__4173));
    ClkMux I__935 (
            .O(N__4244),
            .I(N__4173));
    ClkMux I__934 (
            .O(N__4243),
            .I(N__4173));
    ClkMux I__933 (
            .O(N__4242),
            .I(N__4173));
    ClkMux I__932 (
            .O(N__4241),
            .I(N__4173));
    ClkMux I__931 (
            .O(N__4240),
            .I(N__4173));
    ClkMux I__930 (
            .O(N__4239),
            .I(N__4173));
    ClkMux I__929 (
            .O(N__4238),
            .I(N__4173));
    ClkMux I__928 (
            .O(N__4237),
            .I(N__4173));
    ClkMux I__927 (
            .O(N__4236),
            .I(N__4173));
    ClkMux I__926 (
            .O(N__4235),
            .I(N__4173));
    ClkMux I__925 (
            .O(N__4234),
            .I(N__4173));
    ClkMux I__924 (
            .O(N__4233),
            .I(N__4173));
    ClkMux I__923 (
            .O(N__4232),
            .I(N__4173));
    ClkMux I__922 (
            .O(N__4231),
            .I(N__4173));
    ClkMux I__921 (
            .O(N__4230),
            .I(N__4173));
    GlobalMux I__920 (
            .O(N__4173),
            .I(N__4170));
    gio2CtrlBuf I__919 (
            .O(N__4170),
            .I(i_Clk_c_g));
    IoInMux I__918 (
            .O(N__4167),
            .I(N__4164));
    LocalMux I__917 (
            .O(N__4164),
            .I(N__4161));
    Odrv4 I__916 (
            .O(N__4161),
            .I(r_disp2_i_3));
    InMux I__915 (
            .O(N__4158),
            .I(N__4155));
    LocalMux I__914 (
            .O(N__4155),
            .I(N__4149));
    InMux I__913 (
            .O(N__4154),
            .I(N__4142));
    InMux I__912 (
            .O(N__4153),
            .I(N__4142));
    InMux I__911 (
            .O(N__4152),
            .I(N__4142));
    Span4Mux_v I__910 (
            .O(N__4149),
            .I(N__4135));
    LocalMux I__909 (
            .O(N__4142),
            .I(N__4132));
    InMux I__908 (
            .O(N__4141),
            .I(N__4123));
    InMux I__907 (
            .O(N__4140),
            .I(N__4123));
    InMux I__906 (
            .O(N__4139),
            .I(N__4123));
    InMux I__905 (
            .O(N__4138),
            .I(N__4123));
    Odrv4 I__904 (
            .O(N__4135),
            .I(uart_data_6));
    Odrv4 I__903 (
            .O(N__4132),
            .I(uart_data_6));
    LocalMux I__902 (
            .O(N__4123),
            .I(uart_data_6));
    CascadeMux I__901 (
            .O(N__4116),
            .I(N__4111));
    CascadeMux I__900 (
            .O(N__4115),
            .I(N__4108));
    CascadeMux I__899 (
            .O(N__4114),
            .I(N__4105));
    InMux I__898 (
            .O(N__4111),
            .I(N__4094));
    InMux I__897 (
            .O(N__4108),
            .I(N__4094));
    InMux I__896 (
            .O(N__4105),
            .I(N__4094));
    InMux I__895 (
            .O(N__4104),
            .I(N__4094));
    InMux I__894 (
            .O(N__4103),
            .I(N__4088));
    LocalMux I__893 (
            .O(N__4094),
            .I(N__4085));
    InMux I__892 (
            .O(N__4093),
            .I(N__4078));
    InMux I__891 (
            .O(N__4092),
            .I(N__4078));
    InMux I__890 (
            .O(N__4091),
            .I(N__4078));
    LocalMux I__889 (
            .O(N__4088),
            .I(uart_data_5));
    Odrv12 I__888 (
            .O(N__4085),
            .I(uart_data_5));
    LocalMux I__887 (
            .O(N__4078),
            .I(uart_data_5));
    InMux I__886 (
            .O(N__4071),
            .I(N__4065));
    CascadeMux I__885 (
            .O(N__4070),
            .I(N__4062));
    CascadeMux I__884 (
            .O(N__4069),
            .I(N__4059));
    CascadeMux I__883 (
            .O(N__4068),
            .I(N__4056));
    LocalMux I__882 (
            .O(N__4065),
            .I(N__4052));
    InMux I__881 (
            .O(N__4062),
            .I(N__4045));
    InMux I__880 (
            .O(N__4059),
            .I(N__4045));
    InMux I__879 (
            .O(N__4056),
            .I(N__4045));
    CascadeMux I__878 (
            .O(N__4055),
            .I(N__4039));
    Span4Mux_v I__877 (
            .O(N__4052),
            .I(N__4036));
    LocalMux I__876 (
            .O(N__4045),
            .I(N__4033));
    InMux I__875 (
            .O(N__4044),
            .I(N__4024));
    InMux I__874 (
            .O(N__4043),
            .I(N__4024));
    InMux I__873 (
            .O(N__4042),
            .I(N__4024));
    InMux I__872 (
            .O(N__4039),
            .I(N__4024));
    Odrv4 I__871 (
            .O(N__4036),
            .I(uart_data_7));
    Odrv4 I__870 (
            .O(N__4033),
            .I(uart_data_7));
    LocalMux I__869 (
            .O(N__4024),
            .I(uart_data_7));
    InMux I__868 (
            .O(N__4017),
            .I(N__4014));
    LocalMux I__867 (
            .O(N__4014),
            .I(N__4008));
    InMux I__866 (
            .O(N__4013),
            .I(N__4001));
    InMux I__865 (
            .O(N__4012),
            .I(N__4001));
    InMux I__864 (
            .O(N__4011),
            .I(N__4001));
    Span4Mux_h I__863 (
            .O(N__4008),
            .I(N__3994));
    LocalMux I__862 (
            .O(N__4001),
            .I(N__3991));
    InMux I__861 (
            .O(N__4000),
            .I(N__3982));
    InMux I__860 (
            .O(N__3999),
            .I(N__3982));
    InMux I__859 (
            .O(N__3998),
            .I(N__3982));
    InMux I__858 (
            .O(N__3997),
            .I(N__3982));
    Odrv4 I__857 (
            .O(N__3994),
            .I(uart_data_4));
    Odrv12 I__856 (
            .O(N__3991),
            .I(uart_data_4));
    LocalMux I__855 (
            .O(N__3982),
            .I(uart_data_4));
    IoInMux I__854 (
            .O(N__3975),
            .I(N__3972));
    LocalMux I__853 (
            .O(N__3972),
            .I(N__3969));
    Odrv4 I__852 (
            .O(N__3969),
            .I(r_disp2_i_4));
    InMux I__851 (
            .O(N__3966),
            .I(N__3962));
    CascadeMux I__850 (
            .O(N__3965),
            .I(N__3959));
    LocalMux I__849 (
            .O(N__3962),
            .I(N__3956));
    InMux I__848 (
            .O(N__3959),
            .I(N__3953));
    Odrv4 I__847 (
            .O(N__3956),
            .I(\uart_tx.N_50 ));
    LocalMux I__846 (
            .O(N__3953),
            .I(\uart_tx.N_50 ));
    InMux I__845 (
            .O(N__3948),
            .I(N__3943));
    InMux I__844 (
            .O(N__3947),
            .I(N__3940));
    InMux I__843 (
            .O(N__3946),
            .I(N__3937));
    LocalMux I__842 (
            .O(N__3943),
            .I(\uart_tx.counterZ0Z_0 ));
    LocalMux I__841 (
            .O(N__3940),
            .I(\uart_tx.counterZ0Z_0 ));
    LocalMux I__840 (
            .O(N__3937),
            .I(\uart_tx.counterZ0Z_0 ));
    InMux I__839 (
            .O(N__3930),
            .I(N__3924));
    InMux I__838 (
            .O(N__3929),
            .I(N__3921));
    InMux I__837 (
            .O(N__3928),
            .I(N__3918));
    InMux I__836 (
            .O(N__3927),
            .I(N__3915));
    LocalMux I__835 (
            .O(N__3924),
            .I(\uart_tx.counterZ0Z_1 ));
    LocalMux I__834 (
            .O(N__3921),
            .I(\uart_tx.counterZ0Z_1 ));
    LocalMux I__833 (
            .O(N__3918),
            .I(\uart_tx.counterZ0Z_1 ));
    LocalMux I__832 (
            .O(N__3915),
            .I(\uart_tx.counterZ0Z_1 ));
    InMux I__831 (
            .O(N__3906),
            .I(\uart_tx.un1_counter_5_cry_0 ));
    InMux I__830 (
            .O(N__3903),
            .I(N__3897));
    InMux I__829 (
            .O(N__3902),
            .I(N__3894));
    InMux I__828 (
            .O(N__3901),
            .I(N__3891));
    InMux I__827 (
            .O(N__3900),
            .I(N__3888));
    LocalMux I__826 (
            .O(N__3897),
            .I(\uart_tx.counterZ0Z_2 ));
    LocalMux I__825 (
            .O(N__3894),
            .I(\uart_tx.counterZ0Z_2 ));
    LocalMux I__824 (
            .O(N__3891),
            .I(\uart_tx.counterZ0Z_2 ));
    LocalMux I__823 (
            .O(N__3888),
            .I(\uart_tx.counterZ0Z_2 ));
    InMux I__822 (
            .O(N__3879),
            .I(\uart_tx.un1_counter_5_cry_1 ));
    InMux I__821 (
            .O(N__3876),
            .I(N__3872));
    InMux I__820 (
            .O(N__3875),
            .I(N__3868));
    LocalMux I__819 (
            .O(N__3872),
            .I(N__3865));
    InMux I__818 (
            .O(N__3871),
            .I(N__3862));
    LocalMux I__817 (
            .O(N__3868),
            .I(\uart_tx.counterZ0Z_3 ));
    Odrv4 I__816 (
            .O(N__3865),
            .I(\uart_tx.counterZ0Z_3 ));
    LocalMux I__815 (
            .O(N__3862),
            .I(\uart_tx.counterZ0Z_3 ));
    InMux I__814 (
            .O(N__3855),
            .I(\uart_tx.un1_counter_5_cry_2 ));
    InMux I__813 (
            .O(N__3852),
            .I(N__3846));
    InMux I__812 (
            .O(N__3851),
            .I(N__3841));
    InMux I__811 (
            .O(N__3850),
            .I(N__3841));
    InMux I__810 (
            .O(N__3849),
            .I(N__3838));
    LocalMux I__809 (
            .O(N__3846),
            .I(\uart_tx.counterZ0Z_4 ));
    LocalMux I__808 (
            .O(N__3841),
            .I(\uart_tx.counterZ0Z_4 ));
    LocalMux I__807 (
            .O(N__3838),
            .I(\uart_tx.counterZ0Z_4 ));
    InMux I__806 (
            .O(N__3831),
            .I(\uart_tx.un1_counter_5_cry_3 ));
    InMux I__805 (
            .O(N__3828),
            .I(N__3823));
    InMux I__804 (
            .O(N__3827),
            .I(N__3820));
    InMux I__803 (
            .O(N__3826),
            .I(N__3817));
    LocalMux I__802 (
            .O(N__3823),
            .I(\uart_tx.counterZ0Z_5 ));
    LocalMux I__801 (
            .O(N__3820),
            .I(\uart_tx.counterZ0Z_5 ));
    LocalMux I__800 (
            .O(N__3817),
            .I(\uart_tx.counterZ0Z_5 ));
    InMux I__799 (
            .O(N__3810),
            .I(\uart_tx.un1_counter_5_cry_4 ));
    CascadeMux I__798 (
            .O(N__3807),
            .I(\uart_tx.out_data_2_5_i_m2_ns_1_cascade_ ));
    InMux I__797 (
            .O(N__3804),
            .I(N__3801));
    LocalMux I__796 (
            .O(N__3801),
            .I(\uart_tx.N_57 ));
    InMux I__795 (
            .O(N__3798),
            .I(N__3792));
    InMux I__794 (
            .O(N__3797),
            .I(N__3789));
    InMux I__793 (
            .O(N__3796),
            .I(N__3784));
    InMux I__792 (
            .O(N__3795),
            .I(N__3784));
    LocalMux I__791 (
            .O(N__3792),
            .I(\uart_tx.indexZ0Z_1 ));
    LocalMux I__790 (
            .O(N__3789),
            .I(\uart_tx.indexZ0Z_1 ));
    LocalMux I__789 (
            .O(N__3784),
            .I(\uart_tx.indexZ0Z_1 ));
    CascadeMux I__788 (
            .O(N__3777),
            .I(\uart_tx.N_56_cascade_ ));
    InMux I__787 (
            .O(N__3774),
            .I(N__3769));
    InMux I__786 (
            .O(N__3773),
            .I(N__3765));
    InMux I__785 (
            .O(N__3772),
            .I(N__3762));
    LocalMux I__784 (
            .O(N__3769),
            .I(N__3759));
    InMux I__783 (
            .O(N__3768),
            .I(N__3756));
    LocalMux I__782 (
            .O(N__3765),
            .I(\uart_tx.indexZ0Z_3 ));
    LocalMux I__781 (
            .O(N__3762),
            .I(\uart_tx.indexZ0Z_3 ));
    Odrv12 I__780 (
            .O(N__3759),
            .I(\uart_tx.indexZ0Z_3 ));
    LocalMux I__779 (
            .O(N__3756),
            .I(\uart_tx.indexZ0Z_3 ));
    CascadeMux I__778 (
            .O(N__3747),
            .I(\uart_tx.N_55_cascade_ ));
    InMux I__777 (
            .O(N__3744),
            .I(N__3741));
    LocalMux I__776 (
            .O(N__3741),
            .I(N__3738));
    Span4Mux_h I__775 (
            .O(N__3738),
            .I(N__3735));
    Odrv4 I__774 (
            .O(N__3735),
            .I(\uart_tx.out_data_3_iv_0_a2_1 ));
    IoInMux I__773 (
            .O(N__3732),
            .I(N__3729));
    LocalMux I__772 (
            .O(N__3729),
            .I(N__3726));
    Span4Mux_s3_h I__771 (
            .O(N__3726),
            .I(N__3723));
    Span4Mux_h I__770 (
            .O(N__3723),
            .I(N__3720));
    Odrv4 I__769 (
            .O(N__3720),
            .I(o_UART_TX_c));
    InMux I__768 (
            .O(N__3717),
            .I(N__3714));
    LocalMux I__767 (
            .O(N__3714),
            .I(r_uart_charZ0Z_2));
    InMux I__766 (
            .O(N__3711),
            .I(N__3708));
    LocalMux I__765 (
            .O(N__3708),
            .I(\uart_tx.r_dataZ0Z_2 ));
    InMux I__764 (
            .O(N__3705),
            .I(N__3702));
    LocalMux I__763 (
            .O(N__3702),
            .I(r_uart_charZ0Z_3));
    InMux I__762 (
            .O(N__3699),
            .I(N__3696));
    LocalMux I__761 (
            .O(N__3696),
            .I(\uart_tx.r_dataZ0Z_3 ));
    InMux I__760 (
            .O(N__3693),
            .I(N__3690));
    LocalMux I__759 (
            .O(N__3690),
            .I(r_uart_charZ0Z_6));
    CascadeMux I__758 (
            .O(N__3687),
            .I(N__3684));
    InMux I__757 (
            .O(N__3684),
            .I(N__3681));
    LocalMux I__756 (
            .O(N__3681),
            .I(N__3678));
    Odrv4 I__755 (
            .O(N__3678),
            .I(\uart_tx.r_dataZ0Z_6 ));
    InMux I__754 (
            .O(N__3675),
            .I(N__3672));
    LocalMux I__753 (
            .O(N__3672),
            .I(r_uart_charZ0Z_7));
    InMux I__752 (
            .O(N__3669),
            .I(N__3666));
    LocalMux I__751 (
            .O(N__3666),
            .I(\uart_tx.r_dataZ0Z_7 ));
    CEMux I__750 (
            .O(N__3663),
            .I(N__3660));
    LocalMux I__749 (
            .O(N__3660),
            .I(N__3656));
    CEMux I__748 (
            .O(N__3659),
            .I(N__3652));
    Span4Mux_v I__747 (
            .O(N__3656),
            .I(N__3649));
    CEMux I__746 (
            .O(N__3655),
            .I(N__3646));
    LocalMux I__745 (
            .O(N__3652),
            .I(\uart_tx.r_data_0_sqmuxa ));
    Odrv4 I__744 (
            .O(N__3649),
            .I(\uart_tx.r_data_0_sqmuxa ));
    LocalMux I__743 (
            .O(N__3646),
            .I(\uart_tx.r_data_0_sqmuxa ));
    InMux I__742 (
            .O(N__3639),
            .I(N__3636));
    LocalMux I__741 (
            .O(N__3636),
            .I(N__3633));
    Span4Mux_h I__740 (
            .O(N__3633),
            .I(N__3629));
    InMux I__739 (
            .O(N__3632),
            .I(N__3626));
    Odrv4 I__738 (
            .O(N__3629),
            .I(\uart_rx.r_dataZ0Z_5 ));
    LocalMux I__737 (
            .O(N__3626),
            .I(\uart_rx.r_dataZ0Z_5 ));
    CEMux I__736 (
            .O(N__3621),
            .I(N__3618));
    LocalMux I__735 (
            .O(N__3618),
            .I(N__3613));
    CEMux I__734 (
            .O(N__3617),
            .I(N__3610));
    CEMux I__733 (
            .O(N__3616),
            .I(N__3607));
    Span4Mux_h I__732 (
            .O(N__3613),
            .I(N__3600));
    LocalMux I__731 (
            .O(N__3610),
            .I(N__3600));
    LocalMux I__730 (
            .O(N__3607),
            .I(N__3600));
    Span4Mux_s2_v I__729 (
            .O(N__3600),
            .I(N__3597));
    Odrv4 I__728 (
            .O(N__3597),
            .I(\uart_rx.state_RNIIKQGZ0Z_6 ));
    IoInMux I__727 (
            .O(N__3594),
            .I(N__3591));
    LocalMux I__726 (
            .O(N__3591),
            .I(N__3588));
    Odrv4 I__725 (
            .O(N__3588),
            .I(r_disp2_i_2));
    CascadeMux I__724 (
            .O(N__3585),
            .I(\uart_tx.counter12_7_3_cascade_ ));
    CascadeMux I__723 (
            .O(N__3582),
            .I(N__3579));
    InMux I__722 (
            .O(N__3579),
            .I(N__3573));
    InMux I__721 (
            .O(N__3578),
            .I(N__3573));
    LocalMux I__720 (
            .O(N__3573),
            .I(\uart_tx.counter12_7 ));
    CascadeMux I__719 (
            .O(N__3570),
            .I(\uart_tx.counter12_7_cascade_ ));
    InMux I__718 (
            .O(N__3567),
            .I(N__3564));
    LocalMux I__717 (
            .O(N__3564),
            .I(N__3561));
    Span4Mux_h I__716 (
            .O(N__3561),
            .I(N__3555));
    InMux I__715 (
            .O(N__3560),
            .I(N__3548));
    InMux I__714 (
            .O(N__3559),
            .I(N__3548));
    InMux I__713 (
            .O(N__3558),
            .I(N__3548));
    Odrv4 I__712 (
            .O(N__3555),
            .I(valid_msg));
    LocalMux I__711 (
            .O(N__3548),
            .I(valid_msg));
    CascadeMux I__710 (
            .O(N__3543),
            .I(N__3540));
    InMux I__709 (
            .O(N__3540),
            .I(N__3528));
    InMux I__708 (
            .O(N__3539),
            .I(N__3528));
    InMux I__707 (
            .O(N__3538),
            .I(N__3528));
    InMux I__706 (
            .O(N__3537),
            .I(N__3528));
    LocalMux I__705 (
            .O(N__3528),
            .I(N__3522));
    InMux I__704 (
            .O(N__3527),
            .I(N__3513));
    InMux I__703 (
            .O(N__3526),
            .I(N__3513));
    InMux I__702 (
            .O(N__3525),
            .I(N__3513));
    Span4Mux_v I__701 (
            .O(N__3522),
            .I(N__3510));
    SRMux I__700 (
            .O(N__3521),
            .I(N__3507));
    CascadeMux I__699 (
            .O(N__3520),
            .I(N__3504));
    LocalMux I__698 (
            .O(N__3513),
            .I(N__3500));
    Span4Mux_h I__697 (
            .O(N__3510),
            .I(N__3495));
    LocalMux I__696 (
            .O(N__3507),
            .I(N__3495));
    InMux I__695 (
            .O(N__3504),
            .I(N__3492));
    InMux I__694 (
            .O(N__3503),
            .I(N__3489));
    Span4Mux_h I__693 (
            .O(N__3500),
            .I(N__3481));
    Span4Mux_v I__692 (
            .O(N__3495),
            .I(N__3481));
    LocalMux I__691 (
            .O(N__3492),
            .I(N__3481));
    LocalMux I__690 (
            .O(N__3489),
            .I(N__3478));
    InMux I__689 (
            .O(N__3488),
            .I(N__3475));
    Span4Mux_v I__688 (
            .O(N__3481),
            .I(N__3472));
    Sp12to4 I__687 (
            .O(N__3478),
            .I(N__3466));
    LocalMux I__686 (
            .O(N__3475),
            .I(N__3466));
    Span4Mux_h I__685 (
            .O(N__3472),
            .I(N__3463));
    IoInMux I__684 (
            .O(N__3471),
            .I(N__3460));
    Span12Mux_v I__683 (
            .O(N__3466),
            .I(N__3457));
    IoSpan4Mux I__682 (
            .O(N__3463),
            .I(N__3452));
    LocalMux I__681 (
            .O(N__3460),
            .I(N__3452));
    Odrv12 I__680 (
            .O(N__3457),
            .I(o_LED_1_c));
    Odrv4 I__679 (
            .O(N__3452),
            .I(o_LED_1_c));
    InMux I__678 (
            .O(N__3447),
            .I(N__3442));
    InMux I__677 (
            .O(N__3446),
            .I(N__3439));
    InMux I__676 (
            .O(N__3445),
            .I(N__3436));
    LocalMux I__675 (
            .O(N__3442),
            .I(N__3433));
    LocalMux I__674 (
            .O(N__3439),
            .I(uart_rx_tvalidZ0));
    LocalMux I__673 (
            .O(N__3436),
            .I(uart_rx_tvalidZ0));
    Odrv4 I__672 (
            .O(N__3433),
            .I(uart_rx_tvalidZ0));
    InMux I__671 (
            .O(N__3426),
            .I(N__3422));
    InMux I__670 (
            .O(N__3425),
            .I(N__3416));
    LocalMux I__669 (
            .O(N__3422),
            .I(N__3413));
    InMux I__668 (
            .O(N__3421),
            .I(N__3401));
    InMux I__667 (
            .O(N__3420),
            .I(N__3401));
    InMux I__666 (
            .O(N__3419),
            .I(N__3401));
    LocalMux I__665 (
            .O(N__3416),
            .I(N__3396));
    Span4Mux_h I__664 (
            .O(N__3413),
            .I(N__3396));
    InMux I__663 (
            .O(N__3412),
            .I(N__3385));
    InMux I__662 (
            .O(N__3411),
            .I(N__3385));
    InMux I__661 (
            .O(N__3410),
            .I(N__3385));
    InMux I__660 (
            .O(N__3409),
            .I(N__3385));
    InMux I__659 (
            .O(N__3408),
            .I(N__3385));
    LocalMux I__658 (
            .O(N__3401),
            .I(\uart_tx.stateZ0Z_0 ));
    Odrv4 I__657 (
            .O(N__3396),
            .I(\uart_tx.stateZ0Z_0 ));
    LocalMux I__656 (
            .O(N__3385),
            .I(\uart_tx.stateZ0Z_0 ));
    CascadeMux I__655 (
            .O(N__3378),
            .I(N__3375));
    InMux I__654 (
            .O(N__3375),
            .I(N__3371));
    InMux I__653 (
            .O(N__3374),
            .I(N__3368));
    LocalMux I__652 (
            .O(N__3371),
            .I(\uart_tx.un1_index_ac0_1_0 ));
    LocalMux I__651 (
            .O(N__3368),
            .I(\uart_tx.un1_index_ac0_1_0 ));
    CascadeMux I__650 (
            .O(N__3363),
            .I(N__3355));
    InMux I__649 (
            .O(N__3362),
            .I(N__3352));
    InMux I__648 (
            .O(N__3361),
            .I(N__3349));
    InMux I__647 (
            .O(N__3360),
            .I(N__3346));
    InMux I__646 (
            .O(N__3359),
            .I(N__3343));
    InMux I__645 (
            .O(N__3358),
            .I(N__3338));
    InMux I__644 (
            .O(N__3355),
            .I(N__3338));
    LocalMux I__643 (
            .O(N__3352),
            .I(\uart_tx.indexZ0Z_2 ));
    LocalMux I__642 (
            .O(N__3349),
            .I(\uart_tx.indexZ0Z_2 ));
    LocalMux I__641 (
            .O(N__3346),
            .I(\uart_tx.indexZ0Z_2 ));
    LocalMux I__640 (
            .O(N__3343),
            .I(\uart_tx.indexZ0Z_2 ));
    LocalMux I__639 (
            .O(N__3338),
            .I(\uart_tx.indexZ0Z_2 ));
    InMux I__638 (
            .O(N__3327),
            .I(N__3318));
    InMux I__637 (
            .O(N__3326),
            .I(N__3311));
    InMux I__636 (
            .O(N__3325),
            .I(N__3311));
    InMux I__635 (
            .O(N__3324),
            .I(N__3311));
    InMux I__634 (
            .O(N__3323),
            .I(N__3304));
    InMux I__633 (
            .O(N__3322),
            .I(N__3304));
    InMux I__632 (
            .O(N__3321),
            .I(N__3304));
    LocalMux I__631 (
            .O(N__3318),
            .I(\uart_tx.indexZ0Z_0 ));
    LocalMux I__630 (
            .O(N__3311),
            .I(\uart_tx.indexZ0Z_0 ));
    LocalMux I__629 (
            .O(N__3304),
            .I(\uart_tx.indexZ0Z_0 ));
    InMux I__628 (
            .O(N__3297),
            .I(N__3294));
    LocalMux I__627 (
            .O(N__3294),
            .I(N__3291));
    Span4Mux_h I__626 (
            .O(N__3291),
            .I(N__3288));
    Odrv4 I__625 (
            .O(N__3288),
            .I(\uart_tx.next_state_1_0_m2_i_a2_1_3_0 ));
    CascadeMux I__624 (
            .O(N__3285),
            .I(\uart_tx.next_state_1_0_m2_i_0_0_cascade_ ));
    InMux I__623 (
            .O(N__3282),
            .I(N__3279));
    LocalMux I__622 (
            .O(N__3279),
            .I(\uart_tx.g0_0_3 ));
    CEMux I__621 (
            .O(N__3276),
            .I(N__3273));
    LocalMux I__620 (
            .O(N__3273),
            .I(N__3270));
    Odrv12 I__619 (
            .O(N__3270),
            .I(valid_msg_0));
    IoInMux I__618 (
            .O(N__3267),
            .I(N__3264));
    LocalMux I__617 (
            .O(N__3264),
            .I(N__3261));
    Odrv4 I__616 (
            .O(N__3261),
            .I(r_disp1_i_0));
    IoInMux I__615 (
            .O(N__3258),
            .I(N__3255));
    LocalMux I__614 (
            .O(N__3255),
            .I(N__3252));
    Odrv12 I__613 (
            .O(N__3252),
            .I(r_disp1_i_3));
    InMux I__612 (
            .O(N__3249),
            .I(N__3246));
    LocalMux I__611 (
            .O(N__3246),
            .I(N__3240));
    InMux I__610 (
            .O(N__3245),
            .I(N__3233));
    InMux I__609 (
            .O(N__3244),
            .I(N__3233));
    InMux I__608 (
            .O(N__3243),
            .I(N__3233));
    Span4Mux_h I__607 (
            .O(N__3240),
            .I(N__3226));
    LocalMux I__606 (
            .O(N__3233),
            .I(N__3223));
    InMux I__605 (
            .O(N__3232),
            .I(N__3218));
    InMux I__604 (
            .O(N__3231),
            .I(N__3218));
    InMux I__603 (
            .O(N__3230),
            .I(N__3215));
    InMux I__602 (
            .O(N__3229),
            .I(N__3212));
    Odrv4 I__601 (
            .O(N__3226),
            .I(uart_data_0));
    Odrv12 I__600 (
            .O(N__3223),
            .I(uart_data_0));
    LocalMux I__599 (
            .O(N__3218),
            .I(uart_data_0));
    LocalMux I__598 (
            .O(N__3215),
            .I(uart_data_0));
    LocalMux I__597 (
            .O(N__3212),
            .I(uart_data_0));
    InMux I__596 (
            .O(N__3201),
            .I(N__3198));
    LocalMux I__595 (
            .O(N__3198),
            .I(N__3192));
    InMux I__594 (
            .O(N__3197),
            .I(N__3185));
    InMux I__593 (
            .O(N__3196),
            .I(N__3185));
    InMux I__592 (
            .O(N__3195),
            .I(N__3185));
    Span4Mux_h I__591 (
            .O(N__3192),
            .I(N__3178));
    LocalMux I__590 (
            .O(N__3185),
            .I(N__3175));
    InMux I__589 (
            .O(N__3184),
            .I(N__3170));
    InMux I__588 (
            .O(N__3183),
            .I(N__3170));
    InMux I__587 (
            .O(N__3182),
            .I(N__3167));
    InMux I__586 (
            .O(N__3181),
            .I(N__3164));
    Odrv4 I__585 (
            .O(N__3178),
            .I(uart_data_2));
    Odrv12 I__584 (
            .O(N__3175),
            .I(uart_data_2));
    LocalMux I__583 (
            .O(N__3170),
            .I(uart_data_2));
    LocalMux I__582 (
            .O(N__3167),
            .I(uart_data_2));
    LocalMux I__581 (
            .O(N__3164),
            .I(uart_data_2));
    CascadeMux I__580 (
            .O(N__3153),
            .I(N__3148));
    InMux I__579 (
            .O(N__3152),
            .I(N__3143));
    CascadeMux I__578 (
            .O(N__3151),
            .I(N__3138));
    InMux I__577 (
            .O(N__3148),
            .I(N__3130));
    InMux I__576 (
            .O(N__3147),
            .I(N__3130));
    InMux I__575 (
            .O(N__3146),
            .I(N__3130));
    LocalMux I__574 (
            .O(N__3143),
            .I(N__3127));
    InMux I__573 (
            .O(N__3142),
            .I(N__3124));
    InMux I__572 (
            .O(N__3141),
            .I(N__3121));
    InMux I__571 (
            .O(N__3138),
            .I(N__3116));
    InMux I__570 (
            .O(N__3137),
            .I(N__3116));
    LocalMux I__569 (
            .O(N__3130),
            .I(N__3113));
    Span4Mux_h I__568 (
            .O(N__3127),
            .I(N__3110));
    LocalMux I__567 (
            .O(N__3124),
            .I(uart_data_1));
    LocalMux I__566 (
            .O(N__3121),
            .I(uart_data_1));
    LocalMux I__565 (
            .O(N__3116),
            .I(uart_data_1));
    Odrv4 I__564 (
            .O(N__3113),
            .I(uart_data_1));
    Odrv4 I__563 (
            .O(N__3110),
            .I(uart_data_1));
    CascadeMux I__562 (
            .O(N__3099),
            .I(N__3090));
    CascadeMux I__561 (
            .O(N__3098),
            .I(N__3087));
    InMux I__560 (
            .O(N__3097),
            .I(N__3084));
    CascadeMux I__559 (
            .O(N__3096),
            .I(N__3081));
    CascadeMux I__558 (
            .O(N__3095),
            .I(N__3078));
    CascadeMux I__557 (
            .O(N__3094),
            .I(N__3074));
    InMux I__556 (
            .O(N__3093),
            .I(N__3067));
    InMux I__555 (
            .O(N__3090),
            .I(N__3067));
    InMux I__554 (
            .O(N__3087),
            .I(N__3067));
    LocalMux I__553 (
            .O(N__3084),
            .I(N__3064));
    InMux I__552 (
            .O(N__3081),
            .I(N__3061));
    InMux I__551 (
            .O(N__3078),
            .I(N__3058));
    InMux I__550 (
            .O(N__3077),
            .I(N__3053));
    InMux I__549 (
            .O(N__3074),
            .I(N__3053));
    LocalMux I__548 (
            .O(N__3067),
            .I(N__3050));
    Span4Mux_h I__547 (
            .O(N__3064),
            .I(N__3047));
    LocalMux I__546 (
            .O(N__3061),
            .I(uart_data_3));
    LocalMux I__545 (
            .O(N__3058),
            .I(uart_data_3));
    LocalMux I__544 (
            .O(N__3053),
            .I(uart_data_3));
    Odrv4 I__543 (
            .O(N__3050),
            .I(uart_data_3));
    Odrv4 I__542 (
            .O(N__3047),
            .I(uart_data_3));
    IoInMux I__541 (
            .O(N__3036),
            .I(N__3033));
    LocalMux I__540 (
            .O(N__3033),
            .I(N__3030));
    Odrv4 I__539 (
            .O(N__3030),
            .I(r_disp1_i_2));
    CascadeMux I__538 (
            .O(N__3027),
            .I(\uart_tx.counter12_6_0_cascade_ ));
    InMux I__537 (
            .O(N__3024),
            .I(N__3021));
    LocalMux I__536 (
            .O(N__3021),
            .I(\uart_tx.g0_rn_0 ));
    InMux I__535 (
            .O(N__3018),
            .I(N__3015));
    LocalMux I__534 (
            .O(N__3015),
            .I(\uart_tx.g0_sn ));
    CascadeMux I__533 (
            .O(N__3012),
            .I(N__3009));
    InMux I__532 (
            .O(N__3009),
            .I(N__3006));
    LocalMux I__531 (
            .O(N__3006),
            .I(\uart_tx.r_dataZ0Z_1 ));
    InMux I__530 (
            .O(N__3003),
            .I(N__3000));
    LocalMux I__529 (
            .O(N__3000),
            .I(\uart_tx.r_dataZ0Z_4 ));
    InMux I__528 (
            .O(N__2997),
            .I(N__2994));
    LocalMux I__527 (
            .O(N__2994),
            .I(N__2991));
    Odrv4 I__526 (
            .O(N__2991),
            .I(r_uart_charZ0Z_0));
    InMux I__525 (
            .O(N__2988),
            .I(N__2985));
    LocalMux I__524 (
            .O(N__2985),
            .I(N__2982));
    Odrv12 I__523 (
            .O(N__2982),
            .I(r_uart_charZ0Z_1));
    InMux I__522 (
            .O(N__2979),
            .I(N__2976));
    LocalMux I__521 (
            .O(N__2976),
            .I(N__2973));
    Odrv4 I__520 (
            .O(N__2973),
            .I(r_uart_charZ0Z_4));
    InMux I__519 (
            .O(N__2970),
            .I(N__2967));
    LocalMux I__518 (
            .O(N__2967),
            .I(N__2964));
    Odrv4 I__517 (
            .O(N__2964),
            .I(r_uart_charZ0Z_5));
    InMux I__516 (
            .O(N__2961),
            .I(N__2957));
    CascadeMux I__515 (
            .O(N__2960),
            .I(N__2954));
    LocalMux I__514 (
            .O(N__2957),
            .I(N__2951));
    InMux I__513 (
            .O(N__2954),
            .I(N__2948));
    Span12Mux_s3_v I__512 (
            .O(N__2951),
            .I(N__2945));
    LocalMux I__511 (
            .O(N__2948),
            .I(\uart_rx.r_dataZ0Z_4 ));
    Odrv12 I__510 (
            .O(N__2945),
            .I(\uart_rx.r_dataZ0Z_4 ));
    IoInMux I__509 (
            .O(N__2940),
            .I(N__2937));
    LocalMux I__508 (
            .O(N__2937),
            .I(r_disp1_i_5));
    IoInMux I__507 (
            .O(N__2934),
            .I(N__2931));
    LocalMux I__506 (
            .O(N__2931),
            .I(r_disp1_i_4));
    InMux I__505 (
            .O(N__2928),
            .I(N__2925));
    LocalMux I__504 (
            .O(N__2925),
            .I(CONSTANT_ONE_NET));
    InMux I__503 (
            .O(N__2922),
            .I(N__2919));
    LocalMux I__502 (
            .O(N__2919),
            .I(N__2916));
    Odrv4 I__501 (
            .O(N__2916),
            .I(\uart_tx.r_dataZ0Z_8 ));
    InMux I__500 (
            .O(N__2913),
            .I(N__2910));
    LocalMux I__499 (
            .O(N__2910),
            .I(\uart_tx.r_dataZ0Z_0 ));
    InMux I__498 (
            .O(N__2907),
            .I(N__2904));
    LocalMux I__497 (
            .O(N__2904),
            .I(N__2901));
    Odrv4 I__496 (
            .O(N__2901),
            .I(\uart_tx.r_dataZ0Z_5 ));
    CascadeMux I__495 (
            .O(N__2898),
            .I(\uart_tx.out_data_2_4_i_m2_ns_1_cascade_ ));
    InMux I__494 (
            .O(N__2895),
            .I(N__2889));
    InMux I__493 (
            .O(N__2894),
            .I(N__2886));
    InMux I__492 (
            .O(N__2893),
            .I(N__2881));
    InMux I__491 (
            .O(N__2892),
            .I(N__2881));
    LocalMux I__490 (
            .O(N__2889),
            .I(\uart_rx.timerZ0Z_7 ));
    LocalMux I__489 (
            .O(N__2886),
            .I(\uart_rx.timerZ0Z_7 ));
    LocalMux I__488 (
            .O(N__2881),
            .I(\uart_rx.timerZ0Z_7 ));
    InMux I__487 (
            .O(N__2874),
            .I(\uart_rx.un1_timer_cry_6 ));
    InMux I__486 (
            .O(N__2871),
            .I(bfn_2_13_0_));
    InMux I__485 (
            .O(N__2868),
            .I(N__2864));
    InMux I__484 (
            .O(N__2867),
            .I(N__2861));
    LocalMux I__483 (
            .O(N__2864),
            .I(\uart_rx.timerZ0Z_8 ));
    LocalMux I__482 (
            .O(N__2861),
            .I(\uart_rx.timerZ0Z_8 ));
    SRMux I__481 (
            .O(N__2856),
            .I(N__2852));
    SRMux I__480 (
            .O(N__2855),
            .I(N__2849));
    LocalMux I__479 (
            .O(N__2852),
            .I(N__2846));
    LocalMux I__478 (
            .O(N__2849),
            .I(N__2843));
    Span4Mux_s2_h I__477 (
            .O(N__2846),
            .I(N__2840));
    Odrv4 I__476 (
            .O(N__2843),
            .I(\uart_rx.state_RNIQRIGZ0Z_2 ));
    Odrv4 I__475 (
            .O(N__2840),
            .I(\uart_rx.state_RNIQRIGZ0Z_2 ));
    InMux I__474 (
            .O(N__2835),
            .I(N__2829));
    InMux I__473 (
            .O(N__2834),
            .I(N__2829));
    LocalMux I__472 (
            .O(N__2829),
            .I(N__2825));
    InMux I__471 (
            .O(N__2828),
            .I(N__2822));
    Odrv4 I__470 (
            .O(N__2825),
            .I(\uart_rx.stateZ0Z_6 ));
    LocalMux I__469 (
            .O(N__2822),
            .I(\uart_rx.stateZ0Z_6 ));
    InMux I__468 (
            .O(N__2817),
            .I(N__2812));
    InMux I__467 (
            .O(N__2816),
            .I(N__2809));
    InMux I__466 (
            .O(N__2815),
            .I(N__2806));
    LocalMux I__465 (
            .O(N__2812),
            .I(N__2802));
    LocalMux I__464 (
            .O(N__2809),
            .I(N__2797));
    LocalMux I__463 (
            .O(N__2806),
            .I(N__2797));
    InMux I__462 (
            .O(N__2805),
            .I(N__2794));
    Odrv4 I__461 (
            .O(N__2802),
            .I(\uart_rx.stateZ0Z_0 ));
    Odrv4 I__460 (
            .O(N__2797),
            .I(\uart_rx.stateZ0Z_0 ));
    LocalMux I__459 (
            .O(N__2794),
            .I(\uart_rx.stateZ0Z_0 ));
    InMux I__458 (
            .O(N__2787),
            .I(N__2784));
    LocalMux I__457 (
            .O(N__2784),
            .I(N__2781));
    Span4Mux_s3_v I__456 (
            .O(N__2781),
            .I(N__2777));
    InMux I__455 (
            .O(N__2780),
            .I(N__2774));
    Odrv4 I__454 (
            .O(N__2777),
            .I(\uart_rx.r_dataZ0Z_7 ));
    LocalMux I__453 (
            .O(N__2774),
            .I(\uart_rx.r_dataZ0Z_7 ));
    InMux I__452 (
            .O(N__2769),
            .I(N__2766));
    LocalMux I__451 (
            .O(N__2766),
            .I(N__2762));
    InMux I__450 (
            .O(N__2765),
            .I(N__2759));
    Odrv12 I__449 (
            .O(N__2762),
            .I(\uart_rx.r_dataZ0Z_6 ));
    LocalMux I__448 (
            .O(N__2759),
            .I(\uart_rx.r_dataZ0Z_6 ));
    InMux I__447 (
            .O(N__2754),
            .I(N__2751));
    LocalMux I__446 (
            .O(N__2751),
            .I(N__2747));
    InMux I__445 (
            .O(N__2750),
            .I(N__2744));
    Odrv12 I__444 (
            .O(N__2747),
            .I(\uart_rx.r_dataZ1Z_1 ));
    LocalMux I__443 (
            .O(N__2744),
            .I(\uart_rx.r_dataZ1Z_1 ));
    CascadeMux I__442 (
            .O(N__2739),
            .I(N__2735));
    InMux I__441 (
            .O(N__2738),
            .I(N__2732));
    InMux I__440 (
            .O(N__2735),
            .I(N__2729));
    LocalMux I__439 (
            .O(N__2732),
            .I(N__2726));
    LocalMux I__438 (
            .O(N__2729),
            .I(\uart_rx.r_dataZ0Z_3 ));
    Odrv12 I__437 (
            .O(N__2726),
            .I(\uart_rx.r_dataZ0Z_3 ));
    CascadeMux I__436 (
            .O(N__2721),
            .I(N__2717));
    InMux I__435 (
            .O(N__2720),
            .I(N__2713));
    InMux I__434 (
            .O(N__2717),
            .I(N__2710));
    InMux I__433 (
            .O(N__2716),
            .I(N__2707));
    LocalMux I__432 (
            .O(N__2713),
            .I(\uart_rx.stateZ0Z_2 ));
    LocalMux I__431 (
            .O(N__2710),
            .I(\uart_rx.stateZ0Z_2 ));
    LocalMux I__430 (
            .O(N__2707),
            .I(\uart_rx.stateZ0Z_2 ));
    CascadeMux I__429 (
            .O(N__2700),
            .I(N__2696));
    InMux I__428 (
            .O(N__2699),
            .I(N__2693));
    InMux I__427 (
            .O(N__2696),
            .I(N__2690));
    LocalMux I__426 (
            .O(N__2693),
            .I(\uart_rx.N_123_i ));
    LocalMux I__425 (
            .O(N__2690),
            .I(\uart_rx.N_123_i ));
    InMux I__424 (
            .O(N__2685),
            .I(N__2680));
    InMux I__423 (
            .O(N__2684),
            .I(N__2675));
    InMux I__422 (
            .O(N__2683),
            .I(N__2675));
    LocalMux I__421 (
            .O(N__2680),
            .I(\uart_rx.timerZ0Z_0 ));
    LocalMux I__420 (
            .O(N__2675),
            .I(\uart_rx.timerZ0Z_0 ));
    InMux I__419 (
            .O(N__2670),
            .I(N__2665));
    InMux I__418 (
            .O(N__2669),
            .I(N__2660));
    InMux I__417 (
            .O(N__2668),
            .I(N__2660));
    LocalMux I__416 (
            .O(N__2665),
            .I(\uart_rx.timerZ0Z_1 ));
    LocalMux I__415 (
            .O(N__2660),
            .I(\uart_rx.timerZ0Z_1 ));
    InMux I__414 (
            .O(N__2655),
            .I(\uart_rx.un1_timer_cry_0 ));
    InMux I__413 (
            .O(N__2652),
            .I(N__2646));
    InMux I__412 (
            .O(N__2651),
            .I(N__2643));
    InMux I__411 (
            .O(N__2650),
            .I(N__2638));
    InMux I__410 (
            .O(N__2649),
            .I(N__2638));
    LocalMux I__409 (
            .O(N__2646),
            .I(\uart_rx.timerZ0Z_2 ));
    LocalMux I__408 (
            .O(N__2643),
            .I(\uart_rx.timerZ0Z_2 ));
    LocalMux I__407 (
            .O(N__2638),
            .I(\uart_rx.timerZ0Z_2 ));
    InMux I__406 (
            .O(N__2631),
            .I(\uart_rx.un1_timer_cry_1 ));
    InMux I__405 (
            .O(N__2628),
            .I(N__2623));
    InMux I__404 (
            .O(N__2627),
            .I(N__2620));
    InMux I__403 (
            .O(N__2626),
            .I(N__2617));
    LocalMux I__402 (
            .O(N__2623),
            .I(\uart_rx.timerZ0Z_3 ));
    LocalMux I__401 (
            .O(N__2620),
            .I(\uart_rx.timerZ0Z_3 ));
    LocalMux I__400 (
            .O(N__2617),
            .I(\uart_rx.timerZ0Z_3 ));
    InMux I__399 (
            .O(N__2610),
            .I(\uart_rx.un1_timer_cry_2 ));
    InMux I__398 (
            .O(N__2607),
            .I(N__2600));
    InMux I__397 (
            .O(N__2606),
            .I(N__2595));
    InMux I__396 (
            .O(N__2605),
            .I(N__2595));
    InMux I__395 (
            .O(N__2604),
            .I(N__2592));
    InMux I__394 (
            .O(N__2603),
            .I(N__2589));
    LocalMux I__393 (
            .O(N__2600),
            .I(\uart_rx.timerZ0Z_4 ));
    LocalMux I__392 (
            .O(N__2595),
            .I(\uart_rx.timerZ0Z_4 ));
    LocalMux I__391 (
            .O(N__2592),
            .I(\uart_rx.timerZ0Z_4 ));
    LocalMux I__390 (
            .O(N__2589),
            .I(\uart_rx.timerZ0Z_4 ));
    InMux I__389 (
            .O(N__2580),
            .I(\uart_rx.un1_timer_cry_3 ));
    CascadeMux I__388 (
            .O(N__2577),
            .I(N__2570));
    InMux I__387 (
            .O(N__2576),
            .I(N__2567));
    InMux I__386 (
            .O(N__2575),
            .I(N__2564));
    InMux I__385 (
            .O(N__2574),
            .I(N__2561));
    InMux I__384 (
            .O(N__2573),
            .I(N__2558));
    InMux I__383 (
            .O(N__2570),
            .I(N__2555));
    LocalMux I__382 (
            .O(N__2567),
            .I(\uart_rx.timerZ0Z_5 ));
    LocalMux I__381 (
            .O(N__2564),
            .I(\uart_rx.timerZ0Z_5 ));
    LocalMux I__380 (
            .O(N__2561),
            .I(\uart_rx.timerZ0Z_5 ));
    LocalMux I__379 (
            .O(N__2558),
            .I(\uart_rx.timerZ0Z_5 ));
    LocalMux I__378 (
            .O(N__2555),
            .I(\uart_rx.timerZ0Z_5 ));
    InMux I__377 (
            .O(N__2544),
            .I(\uart_rx.un1_timer_cry_4 ));
    InMux I__376 (
            .O(N__2541),
            .I(N__2537));
    InMux I__375 (
            .O(N__2540),
            .I(N__2534));
    LocalMux I__374 (
            .O(N__2537),
            .I(\uart_rx.timerZ0Z_6 ));
    LocalMux I__373 (
            .O(N__2534),
            .I(\uart_rx.timerZ0Z_6 ));
    InMux I__372 (
            .O(N__2529),
            .I(\uart_rx.un1_timer_cry_5 ));
    InMux I__371 (
            .O(N__2526),
            .I(N__2520));
    InMux I__370 (
            .O(N__2525),
            .I(N__2517));
    InMux I__369 (
            .O(N__2524),
            .I(N__2514));
    InMux I__368 (
            .O(N__2523),
            .I(N__2511));
    LocalMux I__367 (
            .O(N__2520),
            .I(\uart_rx.indexZ0Z_3 ));
    LocalMux I__366 (
            .O(N__2517),
            .I(\uart_rx.indexZ0Z_3 ));
    LocalMux I__365 (
            .O(N__2514),
            .I(\uart_rx.indexZ0Z_3 ));
    LocalMux I__364 (
            .O(N__2511),
            .I(\uart_rx.indexZ0Z_3 ));
    InMux I__363 (
            .O(N__2502),
            .I(N__2496));
    InMux I__362 (
            .O(N__2501),
            .I(N__2493));
    InMux I__361 (
            .O(N__2500),
            .I(N__2490));
    InMux I__360 (
            .O(N__2499),
            .I(N__2487));
    LocalMux I__359 (
            .O(N__2496),
            .I(\uart_rx.indexZ0Z_1 ));
    LocalMux I__358 (
            .O(N__2493),
            .I(\uart_rx.indexZ0Z_1 ));
    LocalMux I__357 (
            .O(N__2490),
            .I(\uart_rx.indexZ0Z_1 ));
    LocalMux I__356 (
            .O(N__2487),
            .I(\uart_rx.indexZ0Z_1 ));
    CascadeMux I__355 (
            .O(N__2478),
            .I(N__2475));
    InMux I__354 (
            .O(N__2475),
            .I(N__2469));
    InMux I__353 (
            .O(N__2474),
            .I(N__2469));
    LocalMux I__352 (
            .O(N__2469),
            .I(\uart_rx.r_datace_0_6 ));
    CascadeMux I__351 (
            .O(N__2466),
            .I(N__2458));
    InMux I__350 (
            .O(N__2465),
            .I(N__2455));
    InMux I__349 (
            .O(N__2464),
            .I(N__2452));
    InMux I__348 (
            .O(N__2463),
            .I(N__2445));
    InMux I__347 (
            .O(N__2462),
            .I(N__2445));
    InMux I__346 (
            .O(N__2461),
            .I(N__2445));
    InMux I__345 (
            .O(N__2458),
            .I(N__2442));
    LocalMux I__344 (
            .O(N__2455),
            .I(\uart_rx.indexZ0Z_2 ));
    LocalMux I__343 (
            .O(N__2452),
            .I(\uart_rx.indexZ0Z_2 ));
    LocalMux I__342 (
            .O(N__2445),
            .I(\uart_rx.indexZ0Z_2 ));
    LocalMux I__341 (
            .O(N__2442),
            .I(\uart_rx.indexZ0Z_2 ));
    InMux I__340 (
            .O(N__2433),
            .I(N__2425));
    InMux I__339 (
            .O(N__2432),
            .I(N__2418));
    InMux I__338 (
            .O(N__2431),
            .I(N__2418));
    InMux I__337 (
            .O(N__2430),
            .I(N__2418));
    InMux I__336 (
            .O(N__2429),
            .I(N__2415));
    InMux I__335 (
            .O(N__2428),
            .I(N__2412));
    LocalMux I__334 (
            .O(N__2425),
            .I(\uart_rx.indexZ0Z_0 ));
    LocalMux I__333 (
            .O(N__2418),
            .I(\uart_rx.indexZ0Z_0 ));
    LocalMux I__332 (
            .O(N__2415),
            .I(\uart_rx.indexZ0Z_0 ));
    LocalMux I__331 (
            .O(N__2412),
            .I(\uart_rx.indexZ0Z_0 ));
    InMux I__330 (
            .O(N__2403),
            .I(N__2397));
    InMux I__329 (
            .O(N__2402),
            .I(N__2397));
    LocalMux I__328 (
            .O(N__2397),
            .I(\uart_rx.r_datace_0_3 ));
    InMux I__327 (
            .O(N__2394),
            .I(N__2383));
    InMux I__326 (
            .O(N__2393),
            .I(N__2383));
    InMux I__325 (
            .O(N__2392),
            .I(N__2380));
    InMux I__324 (
            .O(N__2391),
            .I(N__2375));
    InMux I__323 (
            .O(N__2390),
            .I(N__2368));
    InMux I__322 (
            .O(N__2389),
            .I(N__2368));
    InMux I__321 (
            .O(N__2388),
            .I(N__2368));
    LocalMux I__320 (
            .O(N__2383),
            .I(N__2363));
    LocalMux I__319 (
            .O(N__2380),
            .I(N__2363));
    InMux I__318 (
            .O(N__2379),
            .I(N__2358));
    InMux I__317 (
            .O(N__2378),
            .I(N__2358));
    LocalMux I__316 (
            .O(N__2375),
            .I(\uart_rx.N_122_i ));
    LocalMux I__315 (
            .O(N__2368),
            .I(\uart_rx.N_122_i ));
    Odrv4 I__314 (
            .O(N__2363),
            .I(\uart_rx.N_122_i ));
    LocalMux I__313 (
            .O(N__2358),
            .I(\uart_rx.N_122_i ));
    InMux I__312 (
            .O(N__2349),
            .I(N__2345));
    InMux I__311 (
            .O(N__2348),
            .I(N__2342));
    LocalMux I__310 (
            .O(N__2345),
            .I(\uart_rx.N_147 ));
    LocalMux I__309 (
            .O(N__2342),
            .I(\uart_rx.N_147 ));
    InMux I__308 (
            .O(N__2337),
            .I(N__2331));
    InMux I__307 (
            .O(N__2336),
            .I(N__2326));
    InMux I__306 (
            .O(N__2335),
            .I(N__2326));
    InMux I__305 (
            .O(N__2334),
            .I(N__2323));
    LocalMux I__304 (
            .O(N__2331),
            .I(\uart_rx.N_142 ));
    LocalMux I__303 (
            .O(N__2326),
            .I(\uart_rx.N_142 ));
    LocalMux I__302 (
            .O(N__2323),
            .I(\uart_rx.N_142 ));
    CascadeMux I__301 (
            .O(N__2316),
            .I(N__2309));
    CascadeMux I__300 (
            .O(N__2315),
            .I(N__2305));
    InMux I__299 (
            .O(N__2314),
            .I(N__2299));
    InMux I__298 (
            .O(N__2313),
            .I(N__2292));
    InMux I__297 (
            .O(N__2312),
            .I(N__2292));
    InMux I__296 (
            .O(N__2309),
            .I(N__2292));
    InMux I__295 (
            .O(N__2308),
            .I(N__2287));
    InMux I__294 (
            .O(N__2305),
            .I(N__2287));
    InMux I__293 (
            .O(N__2304),
            .I(N__2284));
    CascadeMux I__292 (
            .O(N__2303),
            .I(N__2281));
    CascadeMux I__291 (
            .O(N__2302),
            .I(N__2278));
    LocalMux I__290 (
            .O(N__2299),
            .I(N__2270));
    LocalMux I__289 (
            .O(N__2292),
            .I(N__2270));
    LocalMux I__288 (
            .O(N__2287),
            .I(N__2270));
    LocalMux I__287 (
            .O(N__2284),
            .I(N__2267));
    InMux I__286 (
            .O(N__2281),
            .I(N__2262));
    InMux I__285 (
            .O(N__2278),
            .I(N__2262));
    CascadeMux I__284 (
            .O(N__2277),
            .I(N__2259));
    Span4Mux_v I__283 (
            .O(N__2270),
            .I(N__2251));
    Span4Mux_s1_h I__282 (
            .O(N__2267),
            .I(N__2251));
    LocalMux I__281 (
            .O(N__2262),
            .I(N__2251));
    InMux I__280 (
            .O(N__2259),
            .I(N__2246));
    InMux I__279 (
            .O(N__2258),
            .I(N__2246));
    Span4Mux_h I__278 (
            .O(N__2251),
            .I(N__2241));
    LocalMux I__277 (
            .O(N__2246),
            .I(N__2241));
    Span4Mux_v I__276 (
            .O(N__2241),
            .I(N__2238));
    Span4Mux_h I__275 (
            .O(N__2238),
            .I(N__2235));
    Span4Mux_h I__274 (
            .O(N__2235),
            .I(N__2232));
    Odrv4 I__273 (
            .O(N__2232),
            .I(i_UART_RX_c));
    InMux I__272 (
            .O(N__2229),
            .I(N__2226));
    LocalMux I__271 (
            .O(N__2226),
            .I(\uart_rx.r_datace_0_5 ));
    SRMux I__270 (
            .O(N__2223),
            .I(N__2220));
    LocalMux I__269 (
            .O(N__2220),
            .I(N__2216));
    SRMux I__268 (
            .O(N__2219),
            .I(N__2213));
    Span4Mux_v I__267 (
            .O(N__2216),
            .I(N__2207));
    LocalMux I__266 (
            .O(N__2213),
            .I(N__2207));
    SRMux I__265 (
            .O(N__2212),
            .I(N__2204));
    Span4Mux_v I__264 (
            .O(N__2207),
            .I(N__2199));
    LocalMux I__263 (
            .O(N__2204),
            .I(N__2199));
    Span4Mux_s1_h I__262 (
            .O(N__2199),
            .I(N__2196));
    Odrv4 I__261 (
            .O(N__2196),
            .I(\uart_rx.state_isoZ0Z_0 ));
    IoInMux I__260 (
            .O(N__2193),
            .I(N__2190));
    LocalMux I__259 (
            .O(N__2190),
            .I(r_disp2_i_1));
    IoInMux I__258 (
            .O(N__2187),
            .I(N__2184));
    LocalMux I__257 (
            .O(N__2184),
            .I(r_disp2_i_0));
    IoInMux I__256 (
            .O(N__2181),
            .I(N__2178));
    LocalMux I__255 (
            .O(N__2178),
            .I(r_disp2_i_6));
    IoInMux I__254 (
            .O(N__2175),
            .I(N__2172));
    LocalMux I__253 (
            .O(N__2172),
            .I(r_disp2_i_5));
    IoInMux I__252 (
            .O(N__2169),
            .I(N__2166));
    LocalMux I__251 (
            .O(N__2166),
            .I(N__2163));
    IoSpan4Mux I__250 (
            .O(N__2163),
            .I(N__2160));
    Odrv4 I__249 (
            .O(N__2160),
            .I(r_disp1_i_1));
    InMux I__248 (
            .O(N__2157),
            .I(N__2153));
    CascadeMux I__247 (
            .O(N__2156),
            .I(N__2150));
    LocalMux I__246 (
            .O(N__2153),
            .I(N__2147));
    InMux I__245 (
            .O(N__2150),
            .I(N__2144));
    Span12Mux_s2_v I__244 (
            .O(N__2147),
            .I(N__2141));
    LocalMux I__243 (
            .O(N__2144),
            .I(\uart_rx.r_dataZ1Z_2 ));
    Odrv12 I__242 (
            .O(N__2141),
            .I(\uart_rx.r_dataZ1Z_2 ));
    InMux I__241 (
            .O(N__2136),
            .I(N__2133));
    LocalMux I__240 (
            .O(N__2133),
            .I(N__2129));
    InMux I__239 (
            .O(N__2132),
            .I(N__2126));
    Odrv12 I__238 (
            .O(N__2129),
            .I(\uart_rx.r_dataZ1Z_0 ));
    LocalMux I__237 (
            .O(N__2126),
            .I(\uart_rx.r_dataZ1Z_0 ));
    IoInMux I__236 (
            .O(N__2121),
            .I(N__2118));
    LocalMux I__235 (
            .O(N__2118),
            .I(r_disp1_i_6));
    InMux I__234 (
            .O(N__2115),
            .I(N__2108));
    InMux I__233 (
            .O(N__2114),
            .I(N__2108));
    InMux I__232 (
            .O(N__2113),
            .I(N__2105));
    LocalMux I__231 (
            .O(N__2108),
            .I(\uart_rx.N_139 ));
    LocalMux I__230 (
            .O(N__2105),
            .I(\uart_rx.N_139 ));
    InMux I__229 (
            .O(N__2100),
            .I(N__2097));
    LocalMux I__228 (
            .O(N__2097),
            .I(\uart_rx.N_136 ));
    InMux I__227 (
            .O(N__2094),
            .I(N__2088));
    InMux I__226 (
            .O(N__2093),
            .I(N__2088));
    LocalMux I__225 (
            .O(N__2088),
            .I(\uart_rx.state_nss_0_i_1_0 ));
    InMux I__224 (
            .O(N__2085),
            .I(N__2082));
    LocalMux I__223 (
            .O(N__2082),
            .I(\uart_rx.state_srsts_i_o2_1_1 ));
    CascadeMux I__222 (
            .O(N__2079),
            .I(\uart_rx.state_srsts_i_a2_1_0_1_cascade_ ));
    InMux I__221 (
            .O(N__2076),
            .I(N__2073));
    LocalMux I__220 (
            .O(N__2073),
            .I(\uart_rx.state_srsts_0_a2_0_1_0_2 ));
    CascadeMux I__219 (
            .O(N__2070),
            .I(\uart_rx.N_130_cascade_ ));
    InMux I__218 (
            .O(N__2067),
            .I(N__2060));
    InMux I__217 (
            .O(N__2066),
            .I(N__2060));
    InMux I__216 (
            .O(N__2065),
            .I(N__2057));
    LocalMux I__215 (
            .O(N__2060),
            .I(\uart_rx.N_109_0 ));
    LocalMux I__214 (
            .O(N__2057),
            .I(\uart_rx.N_109_0 ));
    InMux I__213 (
            .O(N__2052),
            .I(N__2042));
    InMux I__212 (
            .O(N__2051),
            .I(N__2042));
    InMux I__211 (
            .O(N__2050),
            .I(N__2042));
    InMux I__210 (
            .O(N__2049),
            .I(N__2039));
    LocalMux I__209 (
            .O(N__2042),
            .I(\uart_rx.stateZ0Z_1 ));
    LocalMux I__208 (
            .O(N__2039),
            .I(\uart_rx.stateZ0Z_1 ));
    InMux I__207 (
            .O(N__2034),
            .I(N__2031));
    LocalMux I__206 (
            .O(N__2031),
            .I(\uart_rx.state_srsts_0_a2_0_1_4 ));
    CascadeMux I__205 (
            .O(N__2028),
            .I(\uart_rx.state_srsts_0_a2_0_1_4_cascade_ ));
    InMux I__204 (
            .O(N__2025),
            .I(N__2019));
    InMux I__203 (
            .O(N__2024),
            .I(N__2019));
    LocalMux I__202 (
            .O(N__2019),
            .I(N__2015));
    InMux I__201 (
            .O(N__2018),
            .I(N__2012));
    Odrv4 I__200 (
            .O(N__2015),
            .I(\uart_rx.timer_RNIUELTZ0Z_0 ));
    LocalMux I__199 (
            .O(N__2012),
            .I(\uart_rx.timer_RNIUELTZ0Z_0 ));
    CascadeMux I__198 (
            .O(N__2007),
            .I(\uart_rx.N_147_cascade_ ));
    InMux I__197 (
            .O(N__2004),
            .I(N__1998));
    InMux I__196 (
            .O(N__2003),
            .I(N__1998));
    LocalMux I__195 (
            .O(N__1998),
            .I(\uart_rx.state_srsts_0_a2_1_4 ));
    CascadeMux I__194 (
            .O(N__1995),
            .I(\uart_rx.N_136_cascade_ ));
    InMux I__193 (
            .O(N__1992),
            .I(N__1987));
    CascadeMux I__192 (
            .O(N__1991),
            .I(N__1984));
    InMux I__191 (
            .O(N__1990),
            .I(N__1980));
    LocalMux I__190 (
            .O(N__1987),
            .I(N__1977));
    InMux I__189 (
            .O(N__1984),
            .I(N__1974));
    InMux I__188 (
            .O(N__1983),
            .I(N__1971));
    LocalMux I__187 (
            .O(N__1980),
            .I(\uart_rx.stateZ0Z_5 ));
    Odrv12 I__186 (
            .O(N__1977),
            .I(\uart_rx.stateZ0Z_5 ));
    LocalMux I__185 (
            .O(N__1974),
            .I(\uart_rx.stateZ0Z_5 ));
    LocalMux I__184 (
            .O(N__1971),
            .I(\uart_rx.stateZ0Z_5 ));
    CascadeMux I__183 (
            .O(N__1962),
            .I(\uart_rx.state_srsts_0_a2_0_2_2_cascade_ ));
    InMux I__182 (
            .O(N__1959),
            .I(N__1951));
    InMux I__181 (
            .O(N__1958),
            .I(N__1951));
    InMux I__180 (
            .O(N__1957),
            .I(N__1946));
    InMux I__179 (
            .O(N__1956),
            .I(N__1946));
    LocalMux I__178 (
            .O(N__1951),
            .I(\uart_rx.stateZ0Z_3 ));
    LocalMux I__177 (
            .O(N__1946),
            .I(\uart_rx.stateZ0Z_3 ));
    InMux I__176 (
            .O(N__1941),
            .I(\uart_rx.un1_index_cry_2 ));
    InMux I__175 (
            .O(N__1938),
            .I(N__1932));
    InMux I__174 (
            .O(N__1937),
            .I(N__1932));
    LocalMux I__173 (
            .O(N__1932),
            .I(\uart_rx.r_datace_0_2 ));
    CascadeMux I__172 (
            .O(N__1929),
            .I(\uart_rx.N_146_cascade_ ));
    InMux I__171 (
            .O(N__1926),
            .I(N__1923));
    LocalMux I__170 (
            .O(N__1923),
            .I(\uart_rx.N_146 ));
    CascadeMux I__169 (
            .O(N__1920),
            .I(\uart_rx.state_srsts_i_a2_3_3_cascade_ ));
    CascadeMux I__168 (
            .O(N__1917),
            .I(N__1914));
    InMux I__167 (
            .O(N__1914),
            .I(N__1911));
    LocalMux I__166 (
            .O(N__1911),
            .I(\uart_rx.state_srsts_0_a2_2_4 ));
    InMux I__165 (
            .O(N__1908),
            .I(\uart_rx.un1_index_cry_0 ));
    InMux I__164 (
            .O(N__1905),
            .I(\uart_rx.un1_index_cry_1 ));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(\uart_tx.un1_counter_5_cry_7 ),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\uart_rx.un1_timer_cry_7 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uart_rx.index_RNI8GO31_1_0_LC_1_9_2 .C_ON=1'b0;
    defparam \uart_rx.index_RNI8GO31_1_0_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx.index_RNI8GO31_1_0_LC_1_9_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_rx.index_RNI8GO31_1_0_LC_1_9_2  (
            .in0(N__2464),
            .in1(N__2392),
            .in2(_gnd_net_),
            .in3(N__2433),
            .lcout(\uart_rx.r_datace_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.index_RNIA1FR_3_LC_1_9_6 .C_ON=1'b0;
    defparam \uart_rx.index_RNIA1FR_3_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx.index_RNIA1FR_3_LC_1_9_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uart_rx.index_RNIA1FR_3_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(N__2500),
            .in2(_gnd_net_),
            .in3(N__2524),
            .lcout(\uart_rx.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.index_0_LC_1_10_0 .C_ON=1'b1;
    defparam \uart_rx.index_0_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx.index_0_LC_1_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.index_0_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__2429),
            .in2(N__1991),
            .in3(N__1990),
            .lcout(\uart_rx.indexZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\uart_rx.un1_index_cry_0 ),
            .clk(N__4230),
            .ce(),
            .sr(N__2212));
    defparam \uart_rx.index_1_LC_1_10_1 .C_ON=1'b1;
    defparam \uart_rx.index_1_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx.index_1_LC_1_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.index_1_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__2502),
            .in2(_gnd_net_),
            .in3(N__1908),
            .lcout(\uart_rx.indexZ0Z_1 ),
            .ltout(),
            .carryin(\uart_rx.un1_index_cry_0 ),
            .carryout(\uart_rx.un1_index_cry_1 ),
            .clk(N__4230),
            .ce(),
            .sr(N__2212));
    defparam \uart_rx.index_2_LC_1_10_2 .C_ON=1'b1;
    defparam \uart_rx.index_2_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.index_2_LC_1_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.index_2_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__2465),
            .in2(_gnd_net_),
            .in3(N__1905),
            .lcout(\uart_rx.indexZ0Z_2 ),
            .ltout(),
            .carryin(\uart_rx.un1_index_cry_1 ),
            .carryout(\uart_rx.un1_index_cry_2 ),
            .clk(N__4230),
            .ce(),
            .sr(N__2212));
    defparam \uart_rx.index_3_LC_1_10_3 .C_ON=1'b0;
    defparam \uart_rx.index_3_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx.index_3_LC_1_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_rx.index_3_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__2526),
            .in2(_gnd_net_),
            .in3(N__1941),
            .lcout(\uart_rx.indexZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4230),
            .ce(),
            .sr(N__2212));
    defparam \uart_rx.r_data_2_LC_1_10_4 .C_ON=1'b0;
    defparam \uart_rx.r_data_2_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_data_2_LC_1_10_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \uart_rx.r_data_2_LC_1_10_4  (
            .in0(N__1938),
            .in1(N__2308),
            .in2(N__2156),
            .in3(N__2113),
            .lcout(\uart_rx.r_dataZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4230),
            .ce(),
            .sr(N__2212));
    defparam \uart_rx.r_data_0_LC_1_10_5 .C_ON=1'b0;
    defparam \uart_rx.r_data_0_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_data_0_LC_1_10_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \uart_rx.r_data_0_LC_1_10_5  (
            .in0(N__2132),
            .in1(N__1937),
            .in2(N__2315),
            .in3(N__2334),
            .lcout(\uart_rx.r_dataZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4230),
            .ce(),
            .sr(N__2212));
    defparam \uart_rx.state_RNO_0_4_LC_1_11_0 .C_ON=1'b0;
    defparam \uart_rx.state_RNO_0_4_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNO_0_4_LC_1_11_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_rx.state_RNO_0_4_LC_1_11_0  (
            .in0(N__1959),
            .in1(N__2574),
            .in2(_gnd_net_),
            .in3(N__2605),
            .lcout(\uart_rx.state_srsts_0_a2_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNITUIG_2_LC_1_11_1 .C_ON=1'b0;
    defparam \uart_rx.state_RNITUIG_2_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNITUIG_2_LC_1_11_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_rx.state_RNITUIG_2_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__2716),
            .in2(_gnd_net_),
            .in3(N__1958),
            .lcout(\uart_rx.N_146 ),
            .ltout(\uart_rx.N_146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNIGJ841_5_LC_1_11_2 .C_ON=1'b0;
    defparam \uart_rx.state_RNIGJ841_5_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNIGJ841_5_LC_1_11_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uart_rx.state_RNIGJ841_5_LC_1_11_2  (
            .in0(N__2304),
            .in1(N__1983),
            .in2(N__1929),
            .in3(N__2393),
            .lcout(\uart_rx.state_nss_0_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNO_0_3_LC_1_11_3 .C_ON=1'b0;
    defparam \uart_rx.state_RNO_0_3_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNO_0_3_LC_1_11_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \uart_rx.state_RNO_0_3_LC_1_11_3  (
            .in0(N__2606),
            .in1(N__2003),
            .in2(N__2721),
            .in3(N__2576),
            .lcout(),
            .ltout(\uart_rx.state_srsts_i_a2_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_3_LC_1_11_4 .C_ON=1'b0;
    defparam \uart_rx.state_3_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.state_3_LC_1_11_4 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \uart_rx.state_3_LC_1_11_4  (
            .in0(N__3525),
            .in1(N__1926),
            .in2(N__1920),
            .in3(N__2024),
            .lcout(\uart_rx.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4232),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_4_LC_1_11_5 .C_ON=1'b0;
    defparam \uart_rx.state_4_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.state_4_LC_1_11_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uart_rx.state_4_LC_1_11_5  (
            .in0(N__2025),
            .in1(N__2004),
            .in2(N__1917),
            .in3(N__3526),
            .lcout(\uart_rx.N_122_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4232),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.index_RNII0UM1_3_LC_1_11_6 .C_ON=1'b0;
    defparam \uart_rx.index_RNII0UM1_3_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx.index_RNII0UM1_3_LC_1_11_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uart_rx.index_RNII0UM1_3_LC_1_11_6  (
            .in0(N__2525),
            .in1(N__2501),
            .in2(N__2466),
            .in3(N__2428),
            .lcout(\uart_rx.N_147 ),
            .ltout(\uart_rx.N_147_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_5_LC_1_11_7 .C_ON=1'b0;
    defparam \uart_rx.state_5_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx.state_5_LC_1_11_7 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart_rx.state_5_LC_1_11_7  (
            .in0(N__2394),
            .in1(_gnd_net_),
            .in2(N__2007),
            .in3(N__3527),
            .lcout(\uart_rx.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4232),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.timer_RNI1RRB_2_LC_1_12_0 .C_ON=1'b0;
    defparam \uart_rx.timer_RNI1RRB_2_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx.timer_RNI1RRB_2_LC_1_12_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uart_rx.timer_RNI1RRB_2_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__2894),
            .in2(_gnd_net_),
            .in3(N__2651),
            .lcout(\uart_rx.state_srsts_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNI1KSO_6_LC_1_12_1 .C_ON=1'b0;
    defparam \uart_rx.state_RNI1KSO_6_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNI1KSO_6_LC_1_12_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_rx.state_RNI1KSO_6_LC_1_12_1  (
            .in0(N__1957),
            .in1(N__2828),
            .in2(_gnd_net_),
            .in3(N__2378),
            .lcout(\uart_rx.N_136 ),
            .ltout(\uart_rx.N_136_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_0_LC_1_12_2 .C_ON=1'b0;
    defparam \uart_rx.state_0_LC_1_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.state_0_LC_1_12_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \uart_rx.state_0_LC_1_12_2  (
            .in0(N__2093),
            .in1(N__3537),
            .in2(N__1995),
            .in3(N__2066),
            .lcout(\uart_rx.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4233),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_6_LC_1_12_3 .C_ON=1'b0;
    defparam \uart_rx.state_6_LC_1_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx.state_6_LC_1_12_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_rx.state_6_LC_1_12_3  (
            .in0(N__3539),
            .in1(N__2379),
            .in2(_gnd_net_),
            .in3(N__2349),
            .lcout(\uart_rx.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4233),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNO_0_2_LC_1_12_4 .C_ON=1'b0;
    defparam \uart_rx.state_RNO_0_2_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNO_0_2_LC_1_12_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_rx.state_RNO_0_2_LC_1_12_4  (
            .in0(N__2076),
            .in1(N__2575),
            .in2(_gnd_net_),
            .in3(N__2607),
            .lcout(),
            .ltout(\uart_rx.state_srsts_0_a2_0_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_2_LC_1_12_5 .C_ON=1'b0;
    defparam \uart_rx.state_2_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.state_2_LC_1_12_5 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \uart_rx.state_2_LC_1_12_5  (
            .in0(N__3538),
            .in1(N__1992),
            .in2(N__1962),
            .in3(N__2018),
            .lcout(\uart_rx.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4233),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNISTIG_1_LC_1_12_6 .C_ON=1'b0;
    defparam \uart_rx.state_RNISTIG_1_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNISTIG_1_LC_1_12_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_rx.state_RNISTIG_1_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__1956),
            .in2(_gnd_net_),
            .in3(N__2049),
            .lcout(\uart_rx.N_123_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_iso_0_LC_1_12_7 .C_ON=1'b0;
    defparam \uart_rx.state_iso_0_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx.state_iso_0_LC_1_12_7 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \uart_rx.state_iso_0_LC_1_12_7  (
            .in0(N__2067),
            .in1(N__2100),
            .in2(N__3543),
            .in3(N__2094),
            .lcout(\uart_rx.state_isoZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4233),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.timer_RNIOEPH_0_LC_1_13_0 .C_ON=1'b0;
    defparam \uart_rx.timer_RNIOEPH_0_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx.timer_RNIOEPH_0_LC_1_13_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_rx.timer_RNIOEPH_0_LC_1_13_0  (
            .in0(N__2683),
            .in1(N__2668),
            .in2(_gnd_net_),
            .in3(N__2626),
            .lcout(\uart_rx.state_srsts_i_o2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.timer_RNI2MNN_2_LC_1_13_1 .C_ON=1'b0;
    defparam \uart_rx.timer_RNI2MNN_2_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx.timer_RNI2MNN_2_LC_1_13_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uart_rx.timer_RNI2MNN_2_LC_1_13_1  (
            .in0(N__2649),
            .in1(N__2892),
            .in2(N__2577),
            .in3(N__2603),
            .lcout(),
            .ltout(\uart_rx.state_srsts_i_a2_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNITIMT1_1_LC_1_13_2 .C_ON=1'b0;
    defparam \uart_rx.state_RNITIMT1_1_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNITIMT1_1_LC_1_13_2 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \uart_rx.state_RNITIMT1_1_LC_1_13_2  (
            .in0(N__2051),
            .in1(N__2085),
            .in2(N__2079),
            .in3(N__2034),
            .lcout(\uart_rx.N_109_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNO_1_2_LC_1_13_3 .C_ON=1'b0;
    defparam \uart_rx.state_RNO_1_2_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNO_1_2_LC_1_13_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uart_rx.state_RNO_1_2_LC_1_13_3  (
            .in0(N__2650),
            .in1(N__2893),
            .in2(N__2277),
            .in3(N__2050),
            .lcout(\uart_rx.state_srsts_0_a2_0_1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_RNO_0_1_LC_1_13_4 .C_ON=1'b0;
    defparam \uart_rx.state_RNO_0_1_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNO_0_1_LC_1_13_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \uart_rx.state_RNO_0_1_LC_1_13_4  (
            .in0(N__2052),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2258),
            .lcout(),
            .ltout(\uart_rx.N_130_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.state_1_LC_1_13_5 .C_ON=1'b0;
    defparam \uart_rx.state_1_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.state_1_LC_1_13_5 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \uart_rx.state_1_LC_1_13_5  (
            .in0(N__3503),
            .in1(N__2817),
            .in2(N__2070),
            .in3(N__2065),
            .lcout(\uart_rx.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4235),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.timer_RNI60SB_8_LC_1_13_6 .C_ON=1'b0;
    defparam \uart_rx.timer_RNI60SB_8_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx.timer_RNI60SB_8_LC_1_13_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_rx.timer_RNI60SB_8_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__2867),
            .in2(_gnd_net_),
            .in3(N__2540),
            .lcout(\uart_rx.state_srsts_0_a2_0_1_4 ),
            .ltout(\uart_rx.state_srsts_0_a2_0_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.timer_RNIUELT_0_LC_1_13_7 .C_ON=1'b0;
    defparam \uart_rx.timer_RNIUELT_0_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx.timer_RNIUELT_0_LC_1_13_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart_rx.timer_RNIUELT_0_LC_1_13_7  (
            .in0(N__2669),
            .in1(N__2684),
            .in2(N__2028),
            .in3(N__2628),
            .lcout(\uart_rx.timer_RNIUELTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp2_i_1_LC_1_14_2 .C_ON=1'b0;
    defparam \seven_seg.r_disp2_i_1_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp2_i_1_LC_1_14_2 .LUT_INIT=16'b0010100000110010;
    LogicCell40 \seven_seg.r_disp2_i_1_LC_1_14_2  (
            .in0(N__3998),
            .in1(N__4042),
            .in2(N__4114),
            .in3(N__4139),
            .lcout(r_disp2_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4238),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp2_i_0_LC_1_14_3 .C_ON=1'b0;
    defparam \seven_seg.r_disp2_i_0_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp2_i_0_LC_1_14_3 .LUT_INIT=16'b0000100100100001;
    LogicCell40 \seven_seg.r_disp2_i_0_LC_1_14_3  (
            .in0(N__4138),
            .in1(N__4104),
            .in2(N__4055),
            .in3(N__3997),
            .lcout(r_disp2_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4238),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp2_i_6_LC_1_14_4 .C_ON=1'b0;
    defparam \seven_seg.r_disp2_i_6_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp2_i_6_LC_1_14_4 .LUT_INIT=16'b0000100110000010;
    LogicCell40 \seven_seg.r_disp2_i_6_LC_1_14_4  (
            .in0(N__4000),
            .in1(N__4044),
            .in2(N__4116),
            .in3(N__4141),
            .lcout(r_disp2_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4238),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp2_i_5_LC_1_14_6 .C_ON=1'b0;
    defparam \seven_seg.r_disp2_i_5_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp2_i_5_LC_1_14_6 .LUT_INIT=16'b1101011010000000;
    LogicCell40 \seven_seg.r_disp2_i_5_LC_1_14_6  (
            .in0(N__3999),
            .in1(N__4043),
            .in2(N__4115),
            .in3(N__4140),
            .lcout(r_disp2_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4238),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp1_i_1_LC_1_14_7 .C_ON=1'b0;
    defparam \seven_seg.r_disp1_i_1_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp1_i_1_LC_1_14_7 .LUT_INIT=16'b0010110100000100;
    LogicCell40 \seven_seg.r_disp1_i_1_LC_1_14_7  (
            .in0(N__3181),
            .in1(N__3141),
            .in2(N__3095),
            .in3(N__3229),
            .lcout(r_disp1_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4238),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.out_data_2_LC_1_15_6 .C_ON=1'b0;
    defparam \uart_rx.out_data_2_LC_1_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx.out_data_2_LC_1_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.out_data_2_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2157),
            .lcout(uart_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4243),
            .ce(N__3617),
            .sr(_gnd_net_));
    defparam \uart_rx.out_data_0_LC_1_15_7 .C_ON=1'b0;
    defparam \uart_rx.out_data_0_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx.out_data_0_LC_1_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.out_data_0_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2136),
            .lcout(uart_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4243),
            .ce(N__3617),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp1_i_6_LC_1_16_0 .C_ON=1'b0;
    defparam \seven_seg.r_disp1_i_6_LC_1_16_0 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp1_i_6_LC_1_16_0 .LUT_INIT=16'b0110000100000010;
    LogicCell40 \seven_seg.r_disp1_i_6_LC_1_16_0  (
            .in0(N__3182),
            .in1(N__3142),
            .in2(N__3096),
            .in3(N__3230),
            .lcout(r_disp1_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4248),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.r_data_3_LC_2_9_2 .C_ON=1'b0;
    defparam \uart_rx.r_data_3_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_data_3_LC_2_9_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \uart_rx.r_data_3_LC_2_9_2  (
            .in0(N__2403),
            .in1(N__2312),
            .in2(N__2739),
            .in3(N__2114),
            .lcout(\uart_rx.r_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4231),
            .ce(),
            .sr(N__2223));
    defparam \uart_rx.r_data_6_LC_2_9_3 .C_ON=1'b0;
    defparam \uart_rx.r_data_6_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_data_6_LC_2_9_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \uart_rx.r_data_6_LC_2_9_3  (
            .in0(N__2115),
            .in1(N__2314),
            .in2(N__2478),
            .in3(N__2765),
            .lcout(\uart_rx.r_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4231),
            .ce(),
            .sr(N__2223));
    defparam \uart_rx.r_data_4_LC_2_9_4 .C_ON=1'b0;
    defparam \uart_rx.r_data_4_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_data_4_LC_2_9_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \uart_rx.r_data_4_LC_2_9_4  (
            .in0(N__2336),
            .in1(N__2313),
            .in2(N__2960),
            .in3(N__2474),
            .lcout(\uart_rx.r_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4231),
            .ce(),
            .sr(N__2223));
    defparam \uart_rx.r_data_1_LC_2_9_7 .C_ON=1'b0;
    defparam \uart_rx.r_data_1_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_data_1_LC_2_9_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \uart_rx.r_data_1_LC_2_9_7  (
            .in0(N__2750),
            .in1(N__2402),
            .in2(N__2316),
            .in3(N__2335),
            .lcout(\uart_rx.r_dataZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4231),
            .ce(),
            .sr(N__2223));
    defparam \uart_rx.r_data_RNO_0_5_LC_2_10_2 .C_ON=1'b0;
    defparam \uart_rx.r_data_RNO_0_5_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx.r_data_RNO_0_5_LC_2_10_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_rx.r_data_RNO_0_5_LC_2_10_2  (
            .in0(N__2463),
            .in1(N__2390),
            .in2(_gnd_net_),
            .in3(N__2432),
            .lcout(\uart_rx.r_datace_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.index_RNIA1FR_0_3_LC_2_10_3 .C_ON=1'b0;
    defparam \uart_rx.index_RNIA1FR_0_3_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx.index_RNIA1FR_0_3_LC_2_10_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_rx.index_RNIA1FR_0_3_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__2523),
            .in2(_gnd_net_),
            .in3(N__2499),
            .lcout(\uart_rx.N_142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.index_RNI8GO31_0_LC_2_10_4 .C_ON=1'b0;
    defparam \uart_rx.index_RNI8GO31_0_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx.index_RNI8GO31_0_LC_2_10_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_rx.index_RNI8GO31_0_LC_2_10_4  (
            .in0(N__2462),
            .in1(N__2389),
            .in2(_gnd_net_),
            .in3(N__2431),
            .lcout(\uart_rx.r_datace_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.index_RNI8GO31_0_0_LC_2_10_6 .C_ON=1'b0;
    defparam \uart_rx.index_RNI8GO31_0_0_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx.index_RNI8GO31_0_0_LC_2_10_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_rx.index_RNI8GO31_0_0_LC_2_10_6  (
            .in0(N__2461),
            .in1(N__2388),
            .in2(_gnd_net_),
            .in3(N__2430),
            .lcout(\uart_rx.r_datace_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.r_data_7_LC_2_11_1 .C_ON=1'b0;
    defparam \uart_rx.r_data_7_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_data_7_LC_2_11_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \uart_rx.r_data_7_LC_2_11_1  (
            .in0(N__2780),
            .in1(N__2391),
            .in2(N__2303),
            .in3(N__2348),
            .lcout(\uart_rx.r_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4234),
            .ce(),
            .sr(N__2219));
    defparam \uart_rx.r_data_5_LC_2_11_3 .C_ON=1'b0;
    defparam \uart_rx.r_data_5_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_data_5_LC_2_11_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \uart_rx.r_data_5_LC_2_11_3  (
            .in0(N__2337),
            .in1(N__3632),
            .in2(N__2302),
            .in3(N__2229),
            .lcout(\uart_rx.r_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4234),
            .ce(),
            .sr(N__2219));
    defparam \uart_rx.state_RNIQRIG_2_LC_2_11_6 .C_ON=1'b0;
    defparam \uart_rx.state_RNIQRIG_2_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNIQRIG_2_LC_2_11_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_rx.state_RNIQRIG_2_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__2805),
            .in2(_gnd_net_),
            .in3(N__2720),
            .lcout(\uart_rx.state_RNIQRIGZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.out_data_RNO_1_LC_2_11_7 .C_ON=1'b0;
    defparam \uart_tx.out_data_RNO_1_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx.out_data_RNO_1_LC_2_11_7 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \uart_tx.out_data_RNO_1_LC_2_11_7  (
            .in0(N__2922),
            .in1(N__3774),
            .in2(_gnd_net_),
            .in3(N__3426),
            .lcout(\uart_tx.out_data_3_iv_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.timer_0_LC_2_12_0 .C_ON=1'b1;
    defparam \uart_rx.timer_0_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_0_LC_2_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.timer_0_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__2685),
            .in2(N__2700),
            .in3(N__2699),
            .lcout(\uart_rx.timerZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\uart_rx.un1_timer_cry_0 ),
            .clk(N__4236),
            .ce(),
            .sr(N__2856));
    defparam \uart_rx.timer_1_LC_2_12_1 .C_ON=1'b1;
    defparam \uart_rx.timer_1_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_1_LC_2_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.timer_1_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__2670),
            .in2(_gnd_net_),
            .in3(N__2655),
            .lcout(\uart_rx.timerZ0Z_1 ),
            .ltout(),
            .carryin(\uart_rx.un1_timer_cry_0 ),
            .carryout(\uart_rx.un1_timer_cry_1 ),
            .clk(N__4236),
            .ce(),
            .sr(N__2856));
    defparam \uart_rx.timer_2_LC_2_12_2 .C_ON=1'b1;
    defparam \uart_rx.timer_2_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_2_LC_2_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.timer_2_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__2652),
            .in2(_gnd_net_),
            .in3(N__2631),
            .lcout(\uart_rx.timerZ0Z_2 ),
            .ltout(),
            .carryin(\uart_rx.un1_timer_cry_1 ),
            .carryout(\uart_rx.un1_timer_cry_2 ),
            .clk(N__4236),
            .ce(),
            .sr(N__2856));
    defparam \uart_rx.timer_3_LC_2_12_3 .C_ON=1'b1;
    defparam \uart_rx.timer_3_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_3_LC_2_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.timer_3_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__2627),
            .in2(_gnd_net_),
            .in3(N__2610),
            .lcout(\uart_rx.timerZ0Z_3 ),
            .ltout(),
            .carryin(\uart_rx.un1_timer_cry_2 ),
            .carryout(\uart_rx.un1_timer_cry_3 ),
            .clk(N__4236),
            .ce(),
            .sr(N__2856));
    defparam \uart_rx.timer_4_LC_2_12_4 .C_ON=1'b1;
    defparam \uart_rx.timer_4_LC_2_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_4_LC_2_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.timer_4_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__2604),
            .in2(_gnd_net_),
            .in3(N__2580),
            .lcout(\uart_rx.timerZ0Z_4 ),
            .ltout(),
            .carryin(\uart_rx.un1_timer_cry_3 ),
            .carryout(\uart_rx.un1_timer_cry_4 ),
            .clk(N__4236),
            .ce(),
            .sr(N__2856));
    defparam \uart_rx.timer_5_LC_2_12_5 .C_ON=1'b1;
    defparam \uart_rx.timer_5_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_5_LC_2_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.timer_5_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__2573),
            .in2(_gnd_net_),
            .in3(N__2544),
            .lcout(\uart_rx.timerZ0Z_5 ),
            .ltout(),
            .carryin(\uart_rx.un1_timer_cry_4 ),
            .carryout(\uart_rx.un1_timer_cry_5 ),
            .clk(N__4236),
            .ce(),
            .sr(N__2856));
    defparam \uart_rx.timer_6_LC_2_12_6 .C_ON=1'b1;
    defparam \uart_rx.timer_6_LC_2_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_6_LC_2_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.timer_6_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__2541),
            .in2(_gnd_net_),
            .in3(N__2529),
            .lcout(\uart_rx.timerZ0Z_6 ),
            .ltout(),
            .carryin(\uart_rx.un1_timer_cry_5 ),
            .carryout(\uart_rx.un1_timer_cry_6 ),
            .clk(N__4236),
            .ce(),
            .sr(N__2856));
    defparam \uart_rx.timer_7_LC_2_12_7 .C_ON=1'b1;
    defparam \uart_rx.timer_7_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_7_LC_2_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_rx.timer_7_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__2895),
            .in2(_gnd_net_),
            .in3(N__2874),
            .lcout(\uart_rx.timerZ0Z_7 ),
            .ltout(),
            .carryin(\uart_rx.un1_timer_cry_6 ),
            .carryout(\uart_rx.un1_timer_cry_7 ),
            .clk(N__4236),
            .ce(),
            .sr(N__2856));
    defparam \uart_rx.timer_8_LC_2_13_0 .C_ON=1'b0;
    defparam \uart_rx.timer_8_LC_2_13_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx.timer_8_LC_2_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_rx.timer_8_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__2868),
            .in2(_gnd_net_),
            .in3(N__2871),
            .lcout(\uart_rx.timerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4239),
            .ce(),
            .sr(N__2855));
    defparam \uart_rx.state_RNIIKQG_6_LC_2_14_0 .C_ON=1'b0;
    defparam \uart_rx.state_RNIIKQG_6_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \uart_rx.state_RNIIKQG_6_LC_2_14_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_rx.state_RNIIKQG_6_LC_2_14_0  (
            .in0(N__3559),
            .in1(N__2815),
            .in2(_gnd_net_),
            .in3(N__2834),
            .lcout(\uart_rx.state_RNIIKQGZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.r_valid_LC_2_14_5 .C_ON=1'b0;
    defparam \uart_rx.r_valid_LC_2_14_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.r_valid_LC_2_14_5 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \uart_rx.r_valid_LC_2_14_5  (
            .in0(N__2835),
            .in1(N__3560),
            .in2(_gnd_net_),
            .in3(N__2816),
            .lcout(valid_msg),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4244),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.r_valid_RNI3IU7_LC_2_14_7 .C_ON=1'b0;
    defparam \uart_rx.r_valid_RNI3IU7_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx.r_valid_RNI3IU7_LC_2_14_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_rx.r_valid_RNI3IU7_LC_2_14_7  (
            .in0(N__3488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3558),
            .lcout(valid_msg_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.out_data_7_LC_2_15_0 .C_ON=1'b0;
    defparam \uart_rx.out_data_7_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx.out_data_7_LC_2_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.out_data_7_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2787),
            .lcout(uart_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4249),
            .ce(N__3616),
            .sr(_gnd_net_));
    defparam \uart_rx.out_data_6_LC_2_15_1 .C_ON=1'b0;
    defparam \uart_rx.out_data_6_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx.out_data_6_LC_2_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.out_data_6_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2769),
            .lcout(uart_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4249),
            .ce(N__3616),
            .sr(_gnd_net_));
    defparam \uart_rx.out_data_1_LC_2_15_2 .C_ON=1'b0;
    defparam \uart_rx.out_data_1_LC_2_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.out_data_1_LC_2_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.out_data_1_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2754),
            .lcout(uart_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4249),
            .ce(N__3616),
            .sr(_gnd_net_));
    defparam \uart_rx.out_data_3_LC_2_15_4 .C_ON=1'b0;
    defparam \uart_rx.out_data_3_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.out_data_3_LC_2_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.out_data_3_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2738),
            .lcout(uart_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4249),
            .ce(N__3616),
            .sr(_gnd_net_));
    defparam \uart_rx.out_data_4_LC_2_15_6 .C_ON=1'b0;
    defparam \uart_rx.out_data_4_LC_2_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx.out_data_4_LC_2_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.out_data_4_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2961),
            .lcout(uart_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4249),
            .ce(N__3616),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp1_i_5_LC_2_16_2 .C_ON=1'b0;
    defparam \seven_seg.r_disp1_i_5_LC_2_16_2 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp1_i_5_LC_2_16_2 .LUT_INIT=16'b1110010001001000;
    LogicCell40 \seven_seg.r_disp1_i_5_LC_2_16_2  (
            .in0(N__3232),
            .in1(N__3184),
            .in2(N__3151),
            .in3(N__3077),
            .lcout(r_disp1_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4252),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp1_i_4_LC_2_16_5 .C_ON=1'b0;
    defparam \seven_seg.r_disp1_i_4_LC_2_16_5 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp1_i_4_LC_2_16_5 .LUT_INIT=16'b1000000010100100;
    LogicCell40 \seven_seg.r_disp1_i_4_LC_2_16_5  (
            .in0(N__3183),
            .in1(N__3137),
            .in2(N__3094),
            .in3(N__3231),
            .lcout(r_disp1_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4252),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_4_10_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_10_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_10_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.r_data_8_LC_4_11_0 .C_ON=1'b0;
    defparam \uart_tx.r_data_8_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_8_LC_4_11_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_tx.r_data_8_LC_4_11_0  (
            .in0(N__2928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_tx.r_dataZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4240),
            .ce(N__3655),
            .sr(_gnd_net_));
    defparam \uart_tx.r_data_5_LC_4_11_4 .C_ON=1'b0;
    defparam \uart_tx.r_data_5_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_5_LC_4_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.r_data_5_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2970),
            .lcout(\uart_tx.r_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4240),
            .ce(N__3655),
            .sr(_gnd_net_));
    defparam \uart_tx.r_data_0_LC_4_11_5 .C_ON=1'b0;
    defparam \uart_tx.r_data_0_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_0_LC_4_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.r_data_0_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2997),
            .lcout(\uart_tx.r_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4240),
            .ce(N__3655),
            .sr(_gnd_net_));
    defparam \uart_tx.out_data_RNO_5_LC_4_12_1 .C_ON=1'b0;
    defparam \uart_tx.out_data_RNO_5_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx.out_data_RNO_5_LC_4_12_1 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \uart_tx.out_data_RNO_5_LC_4_12_1  (
            .in0(N__3359),
            .in1(N__3322),
            .in2(N__3012),
            .in3(N__2913),
            .lcout(),
            .ltout(\uart_tx.out_data_2_4_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.out_data_RNO_3_LC_4_12_2 .C_ON=1'b0;
    defparam \uart_tx.out_data_RNO_3_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.out_data_RNO_3_LC_4_12_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \uart_tx.out_data_RNO_3_LC_4_12_2  (
            .in0(N__3358),
            .in1(N__2907),
            .in2(N__2898),
            .in3(N__3003),
            .lcout(\uart_tx.N_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.r_data_1_LC_4_12_3 .C_ON=1'b0;
    defparam \uart_tx.r_data_1_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_1_LC_4_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.r_data_1_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2988),
            .lcout(\uart_tx.r_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4245),
            .ce(N__3659),
            .sr(_gnd_net_));
    defparam \uart_tx.r_data_4_LC_4_12_4 .C_ON=1'b0;
    defparam \uart_tx.r_data_4_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_4_LC_4_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.r_data_4_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2979),
            .lcout(\uart_tx.r_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4245),
            .ce(N__3659),
            .sr(_gnd_net_));
    defparam \uart_tx.state_RNO_1_0_LC_4_12_6 .C_ON=1'b0;
    defparam \uart_tx.state_RNO_1_0_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.state_RNO_1_0_LC_4_12_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uart_tx.state_RNO_1_0_LC_4_12_6  (
            .in0(N__3321),
            .in1(N__3795),
            .in2(N__3363),
            .in3(N__3768),
            .lcout(\uart_tx.next_state_1_0_m2_i_a2_1_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.index_RNIB641_1_LC_4_12_7 .C_ON=1'b0;
    defparam \uart_tx.index_RNIB641_1_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx.index_RNIB641_1_LC_4_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_tx.index_RNIB641_1_LC_4_12_7  (
            .in0(N__3796),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3323),
            .lcout(\uart_tx.un1_index_ac0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_uart_char_esr_0_LC_4_14_0.C_ON=1'b0;
    defparam r_uart_char_esr_0_LC_4_14_0.SEQ_MODE=4'b1000;
    defparam r_uart_char_esr_0_LC_4_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 r_uart_char_esr_0_LC_4_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3249),
            .lcout(r_uart_charZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4253),
            .ce(N__3276),
            .sr(N__3521));
    defparam r_uart_char_esr_1_LC_4_14_1.C_ON=1'b0;
    defparam r_uart_char_esr_1_LC_4_14_1.SEQ_MODE=4'b1000;
    defparam r_uart_char_esr_1_LC_4_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 r_uart_char_esr_1_LC_4_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3152),
            .lcout(r_uart_charZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4253),
            .ce(N__3276),
            .sr(N__3521));
    defparam r_uart_char_esr_2_LC_4_14_2.C_ON=1'b0;
    defparam r_uart_char_esr_2_LC_4_14_2.SEQ_MODE=4'b1000;
    defparam r_uart_char_esr_2_LC_4_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 r_uart_char_esr_2_LC_4_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3201),
            .lcout(r_uart_charZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4253),
            .ce(N__3276),
            .sr(N__3521));
    defparam r_uart_char_esr_4_LC_4_14_3.C_ON=1'b0;
    defparam r_uart_char_esr_4_LC_4_14_3.SEQ_MODE=4'b1000;
    defparam r_uart_char_esr_4_LC_4_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 r_uart_char_esr_4_LC_4_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4017),
            .lcout(r_uart_charZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4253),
            .ce(N__3276),
            .sr(N__3521));
    defparam r_uart_char_esr_5_LC_4_14_4.C_ON=1'b0;
    defparam r_uart_char_esr_5_LC_4_14_4.SEQ_MODE=4'b1000;
    defparam r_uart_char_esr_5_LC_4_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 r_uart_char_esr_5_LC_4_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4103),
            .lcout(r_uart_charZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4253),
            .ce(N__3276),
            .sr(N__3521));
    defparam r_uart_char_esr_6_LC_4_14_5.C_ON=1'b0;
    defparam r_uart_char_esr_6_LC_4_14_5.SEQ_MODE=4'b1000;
    defparam r_uart_char_esr_6_LC_4_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 r_uart_char_esr_6_LC_4_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4158),
            .lcout(r_uart_charZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4253),
            .ce(N__3276),
            .sr(N__3521));
    defparam r_uart_char_esr_7_LC_4_14_6.C_ON=1'b0;
    defparam r_uart_char_esr_7_LC_4_14_6.SEQ_MODE=4'b1000;
    defparam r_uart_char_esr_7_LC_4_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 r_uart_char_esr_7_LC_4_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4071),
            .lcout(r_uart_charZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4253),
            .ce(N__3276),
            .sr(N__3521));
    defparam r_uart_char_ess_3_LC_4_14_7.C_ON=1'b0;
    defparam r_uart_char_ess_3_LC_4_14_7.SEQ_MODE=4'b1001;
    defparam r_uart_char_ess_3_LC_4_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 r_uart_char_ess_3_LC_4_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3097),
            .lcout(r_uart_charZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4253),
            .ce(N__3276),
            .sr(N__3521));
    defparam \seven_seg.r_disp1_i_0_LC_4_15_1 .C_ON=1'b0;
    defparam \seven_seg.r_disp1_i_0_LC_4_15_1 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp1_i_0_LC_4_15_1 .LUT_INIT=16'b0000100100100001;
    LogicCell40 \seven_seg.r_disp1_i_0_LC_4_15_1  (
            .in0(N__3195),
            .in1(N__3146),
            .in2(N__3098),
            .in3(N__3243),
            .lcout(r_disp1_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4255),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp1_i_3_LC_4_15_3 .C_ON=1'b0;
    defparam \seven_seg.r_disp1_i_3_LC_4_15_3 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp1_i_3_LC_4_15_3 .LUT_INIT=16'b1000100101000010;
    LogicCell40 \seven_seg.r_disp1_i_3_LC_4_15_3  (
            .in0(N__3197),
            .in1(N__3147),
            .in2(N__3099),
            .in3(N__3245),
            .lcout(r_disp1_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4255),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp1_i_2_LC_4_15_4 .C_ON=1'b0;
    defparam \seven_seg.r_disp1_i_2_LC_4_15_4 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp1_i_2_LC_4_15_4 .LUT_INIT=16'b0000001010101110;
    LogicCell40 \seven_seg.r_disp1_i_2_LC_4_15_4  (
            .in0(N__3244),
            .in1(N__3196),
            .in2(N__3153),
            .in3(N__3093),
            .lcout(r_disp1_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4255),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNI5L34_0_9_LC_5_9_0 .C_ON=1'b0;
    defparam \uart_tx.counter_RNI5L34_0_9_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNI5L34_0_9_LC_5_9_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uart_tx.counter_RNI5L34_0_9_LC_5_9_0  (
            .in0(N__3876),
            .in1(N__3827),
            .in2(N__4467),
            .in3(N__3946),
            .lcout(),
            .ltout(\uart_tx.counter12_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNI9DPM1_1_LC_5_9_1 .C_ON=1'b0;
    defparam \uart_tx.counter_RNI9DPM1_1_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNI9DPM1_1_LC_5_9_1 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \uart_tx.counter_RNI9DPM1_1_LC_5_9_1  (
            .in0(N__3018),
            .in1(N__3024),
            .in2(N__3027),
            .in3(N__3282),
            .lcout(\uart_tx.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.state_RNIT28M_0_LC_5_9_2 .C_ON=1'b0;
    defparam \uart_tx.state_RNIT28M_0_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.state_RNIT28M_0_LC_5_9_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_tx.state_RNIT28M_0_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__3408),
            .in2(_gnd_net_),
            .in3(N__4327),
            .lcout(\uart_tx.g0_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNI1V9O_4_LC_5_9_3 .C_ON=1'b0;
    defparam \uart_tx.counter_RNI1V9O_4_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNI1V9O_4_LC_5_9_3 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \uart_tx.counter_RNI1V9O_4_LC_5_9_3  (
            .in0(N__3409),
            .in1(N__3849),
            .in2(N__4352),
            .in3(N__4560),
            .lcout(\uart_tx.g0_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.state_1_LC_5_9_4 .C_ON=1'b0;
    defparam \uart_tx.state_1_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx.state_1_LC_5_9_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uart_tx.state_1_LC_5_9_4  (
            .in0(N__4406),
            .in1(N__4334),
            .in2(N__3582),
            .in3(N__3411),
            .lcout(\uart_tx.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4237),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.state_RNO_0_0_LC_5_9_5 .C_ON=1'b0;
    defparam \uart_tx.state_RNO_0_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx.state_RNO_0_0_LC_5_9_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \uart_tx.state_RNO_0_0_LC_5_9_5  (
            .in0(N__3410),
            .in1(N__3447),
            .in2(N__4353),
            .in3(N__3297),
            .lcout(),
            .ltout(\uart_tx.next_state_1_0_m2_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.state_0_LC_5_9_6 .C_ON=1'b0;
    defparam \uart_tx.state_0_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_tx.state_0_LC_5_9_6 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \uart_tx.state_0_LC_5_9_6  (
            .in0(N__3578),
            .in1(N__4405),
            .in2(N__3285),
            .in3(N__3412),
            .lcout(\uart_tx.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4237),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNI6M34_0_1_LC_5_9_7 .C_ON=1'b0;
    defparam \uart_tx.counter_RNI6M34_0_1_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNI6M34_0_1_LC_5_9_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uart_tx.counter_RNI6M34_0_1_LC_5_9_7  (
            .in0(N__3900),
            .in1(N__3927),
            .in2(N__4531),
            .in3(N__4494),
            .lcout(\uart_tx.g0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNI5L34_9_LC_5_10_0 .C_ON=1'b0;
    defparam \uart_tx.counter_RNI5L34_9_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNI5L34_9_LC_5_10_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uart_tx.counter_RNI5L34_9_LC_5_10_0  (
            .in0(N__3826),
            .in1(N__3871),
            .in2(N__4463),
            .in3(N__3947),
            .lcout(\uart_tx.counter12_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNI1V9O_0_4_LC_5_10_1 .C_ON=1'b0;
    defparam \uart_tx.counter_RNI1V9O_0_4_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNI1V9O_0_4_LC_5_10_1 .LUT_INIT=16'b0000000010110011;
    LogicCell40 \uart_tx.counter_RNI1V9O_0_4_LC_5_10_1  (
            .in0(N__3850),
            .in1(N__4346),
            .in2(N__4571),
            .in3(N__3419),
            .lcout(\uart_tx.counter_RNI1V9O_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.state_RNIT28M_0_0_LC_5_10_2 .C_ON=1'b0;
    defparam \uart_tx.state_RNIT28M_0_0_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.state_RNIT28M_0_0_LC_5_10_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uart_tx.state_RNIT28M_0_0_LC_5_10_2  (
            .in0(N__3421),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4356),
            .lcout(\uart_tx.tready5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNI6M34_1_LC_5_10_3 .C_ON=1'b0;
    defparam \uart_tx.counter_RNI6M34_1_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNI6M34_1_LC_5_10_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uart_tx.counter_RNI6M34_1_LC_5_10_3  (
            .in0(N__3902),
            .in1(N__4496),
            .in2(N__4535),
            .in3(N__3929),
            .lcout(\uart_tx.counter_RNI6M34Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNI6M34_1_1_LC_5_10_4 .C_ON=1'b0;
    defparam \uart_tx.counter_RNI6M34_1_1_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNI6M34_1_1_LC_5_10_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uart_tx.counter_RNI6M34_1_1_LC_5_10_4  (
            .in0(N__3901),
            .in1(N__3928),
            .in2(N__4536),
            .in3(N__4495),
            .lcout(),
            .ltout(\uart_tx.counter12_7_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_RNIAI56_4_LC_5_10_5 .C_ON=1'b0;
    defparam \uart_tx.counter_RNIAI56_4_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx.counter_RNIAI56_4_LC_5_10_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uart_tx.counter_RNIAI56_4_LC_5_10_5  (
            .in0(N__3851),
            .in1(_gnd_net_),
            .in2(N__3585),
            .in3(N__4572),
            .lcout(\uart_tx.counter12_7 ),
            .ltout(\uart_tx.counter12_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.state_RNICAH01_0_LC_5_10_6 .C_ON=1'b0;
    defparam \uart_tx.state_RNICAH01_0_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.state_RNICAH01_0_LC_5_10_6 .LUT_INIT=16'b0111000100010001;
    LogicCell40 \uart_tx.state_RNICAH01_0_LC_5_10_6  (
            .in0(N__3420),
            .in1(N__4355),
            .in2(N__3570),
            .in3(N__4407),
            .lcout(\uart_tx.state_RNICAH01Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam uart_rx_tvalid_LC_5_10_7.C_ON=1'b0;
    defparam uart_rx_tvalid_LC_5_10_7.SEQ_MODE=4'b1000;
    defparam uart_rx_tvalid_LC_5_10_7.LUT_INIT=16'b0000010100001100;
    LogicCell40 uart_rx_tvalid_LC_5_10_7 (
            .in0(N__4269),
            .in1(N__3567),
            .in2(N__3520),
            .in3(N__3446),
            .lcout(uart_rx_tvalidZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4241),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.index_3_LC_5_11_0 .C_ON=1'b0;
    defparam \uart_tx.index_3_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.index_3_LC_5_11_0 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \uart_tx.index_3_LC_5_11_0  (
            .in0(N__4378),
            .in1(N__3773),
            .in2(N__3378),
            .in3(N__3362),
            .lcout(\uart_tx.indexZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4246),
            .ce(),
            .sr(N__4296));
    defparam \uart_tx.index_1_LC_5_11_1 .C_ON=1'b0;
    defparam \uart_tx.index_1_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.index_1_LC_5_11_1 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \uart_tx.index_1_LC_5_11_1  (
            .in0(N__3798),
            .in1(N__4377),
            .in2(_gnd_net_),
            .in3(N__3327),
            .lcout(\uart_tx.indexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4246),
            .ce(),
            .sr(N__4296));
    defparam \uart_tx.state_RNI562Q_0_LC_5_11_2 .C_ON=1'b0;
    defparam \uart_tx.state_RNI562Q_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.state_RNI562Q_0_LC_5_11_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_tx.state_RNI562Q_0_LC_5_11_2  (
            .in0(N__4354),
            .in1(N__3445),
            .in2(_gnd_net_),
            .in3(N__3425),
            .lcout(\uart_tx.r_data_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.index_0_LC_5_12_2 .C_ON=1'b0;
    defparam \uart_tx.index_0_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx.index_0_LC_5_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \uart_tx.index_0_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__4379),
            .in2(_gnd_net_),
            .in3(N__3326),
            .lcout(\uart_tx.indexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4250),
            .ce(),
            .sr(N__4295));
    defparam \uart_tx.index_2_LC_5_12_3 .C_ON=1'b0;
    defparam \uart_tx.index_2_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.index_2_LC_5_12_3 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \uart_tx.index_2_LC_5_12_3  (
            .in0(N__3361),
            .in1(N__3374),
            .in2(_gnd_net_),
            .in3(N__4380),
            .lcout(\uart_tx.indexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4250),
            .ce(),
            .sr(N__4295));
    defparam \uart_tx.out_data_RNO_4_LC_5_12_4 .C_ON=1'b0;
    defparam \uart_tx.out_data_RNO_4_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx.out_data_RNO_4_LC_5_12_4 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \uart_tx.out_data_RNO_4_LC_5_12_4  (
            .in0(N__3360),
            .in1(N__3324),
            .in2(N__3687),
            .in3(N__3711),
            .lcout(),
            .ltout(\uart_tx.out_data_2_5_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.out_data_RNO_2_LC_5_12_5 .C_ON=1'b0;
    defparam \uart_tx.out_data_RNO_2_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx.out_data_RNO_2_LC_5_12_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \uart_tx.out_data_RNO_2_LC_5_12_5  (
            .in0(N__3325),
            .in1(N__3669),
            .in2(N__3807),
            .in3(N__3699),
            .lcout(),
            .ltout(\uart_tx.N_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.out_data_RNO_0_LC_5_12_6 .C_ON=1'b0;
    defparam \uart_tx.out_data_RNO_0_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.out_data_RNO_0_LC_5_12_6 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \uart_tx.out_data_RNO_0_LC_5_12_6  (
            .in0(N__3804),
            .in1(N__3797),
            .in2(N__3777),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\uart_tx.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.out_data_LC_5_12_7 .C_ON=1'b0;
    defparam \uart_tx.out_data_LC_5_12_7 .SEQ_MODE=4'b1001;
    defparam \uart_tx.out_data_LC_5_12_7 .LUT_INIT=16'b0010000010101010;
    LogicCell40 \uart_tx.out_data_LC_5_12_7  (
            .in0(N__4357),
            .in1(N__3772),
            .in2(N__3747),
            .in3(N__3744),
            .lcout(o_UART_TX_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4250),
            .ce(),
            .sr(N__4295));
    defparam \uart_tx.r_data_2_LC_5_13_0 .C_ON=1'b0;
    defparam \uart_tx.r_data_2_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_2_LC_5_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.r_data_2_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3717),
            .lcout(\uart_tx.r_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4254),
            .ce(N__3663),
            .sr(_gnd_net_));
    defparam \uart_tx.r_data_3_LC_5_13_1 .C_ON=1'b0;
    defparam \uart_tx.r_data_3_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_3_LC_5_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.r_data_3_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3705),
            .lcout(\uart_tx.r_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4254),
            .ce(N__3663),
            .sr(_gnd_net_));
    defparam \uart_tx.r_data_6_LC_5_13_2 .C_ON=1'b0;
    defparam \uart_tx.r_data_6_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_6_LC_5_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.r_data_6_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3693),
            .lcout(\uart_tx.r_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4254),
            .ce(N__3663),
            .sr(_gnd_net_));
    defparam \uart_tx.r_data_7_LC_5_13_3 .C_ON=1'b0;
    defparam \uart_tx.r_data_7_LC_5_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.r_data_7_LC_5_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_tx.r_data_7_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3675),
            .lcout(\uart_tx.r_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4254),
            .ce(N__3663),
            .sr(_gnd_net_));
    defparam \uart_rx.out_data_5_LC_5_14_4 .C_ON=1'b0;
    defparam \uart_rx.out_data_5_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.out_data_5_LC_5_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.out_data_5_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3639),
            .lcout(uart_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4256),
            .ce(N__3621),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp2_i_2_LC_5_15_1 .C_ON=1'b0;
    defparam \seven_seg.r_disp2_i_2_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp2_i_2_LC_5_15_1 .LUT_INIT=16'b0001111100000010;
    LogicCell40 \seven_seg.r_disp2_i_2_LC_5_15_1  (
            .in0(N__4152),
            .in1(N__4091),
            .in2(N__4068),
            .in3(N__4011),
            .lcout(r_disp2_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4257),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp2_i_3_LC_5_15_3 .C_ON=1'b0;
    defparam \seven_seg.r_disp2_i_3_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp2_i_3_LC_5_15_3 .LUT_INIT=16'b1000100101000010;
    LogicCell40 \seven_seg.r_disp2_i_3_LC_5_15_3  (
            .in0(N__4153),
            .in1(N__4092),
            .in2(N__4069),
            .in3(N__4012),
            .lcout(r_disp2_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4257),
            .ce(),
            .sr(_gnd_net_));
    defparam \seven_seg.r_disp2_i_4_LC_5_15_7 .C_ON=1'b0;
    defparam \seven_seg.r_disp2_i_4_LC_5_15_7 .SEQ_MODE=4'b1000;
    defparam \seven_seg.r_disp2_i_4_LC_5_15_7 .LUT_INIT=16'b1000000010100100;
    LogicCell40 \seven_seg.r_disp2_i_4_LC_5_15_7  (
            .in0(N__4154),
            .in1(N__4093),
            .in2(N__4070),
            .in3(N__4013),
            .lcout(r_disp2_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4257),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.counter_0_LC_6_9_0 .C_ON=1'b1;
    defparam \uart_tx.counter_0_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_0_LC_6_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_0_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__3948),
            .in2(N__3965),
            .in3(N__3966),
            .lcout(\uart_tx.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\uart_tx.un1_counter_5_cry_0 ),
            .clk(N__4242),
            .ce(),
            .sr(N__4440));
    defparam \uart_tx.counter_1_LC_6_9_1 .C_ON=1'b1;
    defparam \uart_tx.counter_1_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_1_LC_6_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_1_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__3930),
            .in2(_gnd_net_),
            .in3(N__3906),
            .lcout(\uart_tx.counterZ0Z_1 ),
            .ltout(),
            .carryin(\uart_tx.un1_counter_5_cry_0 ),
            .carryout(\uart_tx.un1_counter_5_cry_1 ),
            .clk(N__4242),
            .ce(),
            .sr(N__4440));
    defparam \uart_tx.counter_2_LC_6_9_2 .C_ON=1'b1;
    defparam \uart_tx.counter_2_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_2_LC_6_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_2_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__3903),
            .in2(_gnd_net_),
            .in3(N__3879),
            .lcout(\uart_tx.counterZ0Z_2 ),
            .ltout(),
            .carryin(\uart_tx.un1_counter_5_cry_1 ),
            .carryout(\uart_tx.un1_counter_5_cry_2 ),
            .clk(N__4242),
            .ce(),
            .sr(N__4440));
    defparam \uart_tx.counter_3_LC_6_9_3 .C_ON=1'b1;
    defparam \uart_tx.counter_3_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_3_LC_6_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_3_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__3875),
            .in2(_gnd_net_),
            .in3(N__3855),
            .lcout(\uart_tx.counterZ0Z_3 ),
            .ltout(),
            .carryin(\uart_tx.un1_counter_5_cry_2 ),
            .carryout(\uart_tx.un1_counter_5_cry_3 ),
            .clk(N__4242),
            .ce(),
            .sr(N__4440));
    defparam \uart_tx.counter_4_LC_6_9_4 .C_ON=1'b1;
    defparam \uart_tx.counter_4_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_4_LC_6_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_4_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__3852),
            .in2(_gnd_net_),
            .in3(N__3831),
            .lcout(\uart_tx.counterZ0Z_4 ),
            .ltout(),
            .carryin(\uart_tx.un1_counter_5_cry_3 ),
            .carryout(\uart_tx.un1_counter_5_cry_4 ),
            .clk(N__4242),
            .ce(),
            .sr(N__4440));
    defparam \uart_tx.counter_5_LC_6_9_5 .C_ON=1'b1;
    defparam \uart_tx.counter_5_LC_6_9_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_5_LC_6_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_5_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__3828),
            .in2(_gnd_net_),
            .in3(N__3810),
            .lcout(\uart_tx.counterZ0Z_5 ),
            .ltout(),
            .carryin(\uart_tx.un1_counter_5_cry_4 ),
            .carryout(\uart_tx.un1_counter_5_cry_5 ),
            .clk(N__4242),
            .ce(),
            .sr(N__4440));
    defparam \uart_tx.counter_6_LC_6_9_6 .C_ON=1'b1;
    defparam \uart_tx.counter_6_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_6_LC_6_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_6_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(N__4567),
            .in2(_gnd_net_),
            .in3(N__4539),
            .lcout(\uart_tx.counterZ0Z_6 ),
            .ltout(),
            .carryin(\uart_tx.un1_counter_5_cry_5 ),
            .carryout(\uart_tx.un1_counter_5_cry_6 ),
            .clk(N__4242),
            .ce(),
            .sr(N__4440));
    defparam \uart_tx.counter_7_LC_6_9_7 .C_ON=1'b1;
    defparam \uart_tx.counter_7_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_7_LC_6_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_7_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(N__4530),
            .in2(_gnd_net_),
            .in3(N__4500),
            .lcout(\uart_tx.counterZ0Z_7 ),
            .ltout(),
            .carryin(\uart_tx.un1_counter_5_cry_6 ),
            .carryout(\uart_tx.un1_counter_5_cry_7 ),
            .clk(N__4242),
            .ce(),
            .sr(N__4440));
    defparam \uart_tx.counter_8_LC_6_10_0 .C_ON=1'b1;
    defparam \uart_tx.counter_8_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_8_LC_6_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.counter_8_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__4497),
            .in2(_gnd_net_),
            .in3(N__4473),
            .lcout(\uart_tx.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\uart_tx.un1_counter_5_cry_8 ),
            .clk(N__4247),
            .ce(),
            .sr(N__4436));
    defparam \uart_tx.counter_9_LC_6_10_1 .C_ON=1'b0;
    defparam \uart_tx.counter_9_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.counter_9_LC_6_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_tx.counter_9_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__4462),
            .in2(_gnd_net_),
            .in3(N__4470),
            .lcout(\uart_tx.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4247),
            .ce(),
            .sr(N__4436));
    defparam \uart_tx.state_RNIBCLB1_1_LC_6_11_6 .C_ON=1'b0;
    defparam \uart_tx.state_RNIBCLB1_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.state_RNIBCLB1_1_LC_6_11_6 .LUT_INIT=16'b0100111111001111;
    LogicCell40 \uart_tx.state_RNIBCLB1_1_LC_6_11_6  (
            .in0(N__4422),
            .in1(N__4358),
            .in2(N__4416),
            .in3(N__4401),
            .lcout(\uart_tx.N_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.tready_LC_6_11_7 .C_ON=1'b0;
    defparam \uart_tx.tready_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.tready_LC_6_11_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \uart_tx.tready_LC_6_11_7  (
            .in0(N__4359),
            .in1(N__4268),
            .in2(_gnd_net_),
            .in3(N__4285),
            .lcout(uart_tx_tready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4251),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
